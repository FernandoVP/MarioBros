library ieee;

use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity pipe1_ROM is

	Port(
	
		dir_y : in integer;
		dir_x : in integer;
		
		dat_R : out std_logic_vector( 7 downto 0 );
		dat_G : out std_logic_vector( 7 downto 0 );
		dat_B : out std_logic_vector( 7 downto 0 )
		
	);

end pipe1_ROM;

architecture comp of pipe1_ROM is

	type arreglo is array( 0 to 30 ) of std_logic_vector( 0 to 7 );

	type ROM is array( 0 to 30 ) of arreglo;

	constant pipe_R : ROM :=
	(
	
		(x"08",x"00",x"01",x"00",x"07",x"01",x"02",x"04",x"00",x"05",x"06",x"00",x"0C",x"00",x"02",x"0C",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"00",x"0C",x"06",x"04",x"01",x"04",x"09"),
		(x"07",x"A2",x"AB",x"A5",x"A5",x"A9",x"9A",x"A5",x"B0",x"A0",x"9C",x"AD",x"A2",x"A9",x"A5",x"9D",x"A6",x"A6",x"A6",x"A6",x"A6",x"A6",x"A6",x"A6",x"A5",x"97",x"AF",x"9D",x"AB",x"A8",x"A2"),
		(x"00",x"25",x"14",x"14",x"0E",x"29",x"AB",x"A7",x"9F",x"AC",x"B4",x"A6",x"15",x"16",x"1F",x"1A",x"1B",x"1B",x"1B",x"1B",x"1B",x"1B",x"1B",x"1B",x"23",x"0E",x"17",x"23",x"1C",x"0E",x"1E"),
		(x"01",x"AA",x"B1",x"AC",x"1C",x"1A",x"94",x"9E",x"93",x"A1",x"97",x"94",x"21",x"A6",x"9D",x"21",x"1B",x"1B",x"1B",x"1B",x"1B",x"1B",x"1B",x"1B",x"21",x"A8",x"28",x"A8",x"20",x"97",x"A7"),
		(x"12",x"9F",x"A7",x"9C",x"1E",x"18",x"AC",x"AD",x"9E",x"AB",x"A8",x"AB",x"0E",x"A4",x"A1",x"1B",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1D",x"18",x"92",x"1F",x"9A",x"AA",x"A3"),
		(x"00",x"A0",x"A5",x"9A",x"1F",x"1A",x"9C",x"9D",x"AB",x"A8",x"9F",x"AB",x"16",x"B4",x"AA",x"16",x"1B",x"1B",x"1B",x"1B",x"1B",x"1B",x"1B",x"1B",x"21",x"9D",x"25",x"AE",x"22",x"A8",x"A0"),
		(x"03",x"9E",x"98",x"9C",x"29",x"25",x"A2",x"9D",x"AB",x"9D",x"97",x"AB",x"1E",x"A3",x"9F",x"1E",x"1A",x"1A",x"1A",x"1A",x"1A",x"1A",x"1A",x"1A",x"1F",x"12",x"9B",x"1A",x"AA",x"A4",x"9F"),
		(x"09",x"AA",x"A6",x"9E",x"22",x"11",x"A7",x"AB",x"96",x"AA",x"AF",x"A1",x"15",x"A0",x"A5",x"20",x"1D",x"1D",x"1D",x"1D",x"1D",x"1D",x"1D",x"1D",x"1E",x"9B",x"2A",x"A4",x"0F",x"A0",x"A0"),
		(x"00",x"B3",x"A2",x"A5",x"21",x"12",x"9F",x"A7",x"A6",x"9F",x"A7",x"A3",x"1C",x"9E",x"A4",x"1B",x"1A",x"1A",x"1A",x"1A",x"1A",x"1A",x"1A",x"1A",x"1D",x"0E",x"A0",x"24",x"9A",x"98",x"B0"),
		(x"00",x"9F",x"A7",x"A2",x"23",x"1D",x"99",x"A9",x"9E",x"A7",x"9C",x"A0",x"2C",x"9F",x"96",x"2D",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"1F",x"2B",x"A8",x"26",x"9D",x"32",x"9E",x"B0"),
		(x"0B",x"AC",x"A3",x"9E",x"1D",x"15",x"A8",x"A0",x"A4",x"A6",x"A2",x"AB",x"20",x"A0",x"9D",x"26",x"19",x"19",x"19",x"19",x"19",x"19",x"19",x"19",x"0B",x"13",x"9C",x"18",x"9B",x"A6",x"A0"),
		(x"11",x"98",x"A1",x"9E",x"1A",x"18",x"9E",x"AB",x"A3",x"A3",x"98",x"AD",x"1D",x"A1",x"95",x"29",x"1C",x"1C",x"1C",x"1C",x"1C",x"1C",x"1C",x"1C",x"21",x"AB",x"21",x"A5",x"13",x"A9",x"AE"),
		(x"04",x"9C",x"AF",x"A2",x"1B",x"22",x"9C",x"A4",x"A1",x"AB",x"A5",x"A7",x"12",x"A6",x"9F",x"17",x"1D",x"1D",x"1D",x"1D",x"1D",x"1D",x"1D",x"1D",x"19",x"1C",x"AC",x"1F",x"9F",x"AD",x"A0"),
		(x"00",x"96",x"A9",x"9D",x"2B",x"2E",x"9E",x"AB",x"A1",x"A1",x"A9",x"A1",x"26",x"A1",x"AA",x"26",x"1B",x"1B",x"1B",x"1B",x"1B",x"1B",x"1B",x"1B",x"28",x"9A",x"24",x"9C",x"1C",x"AD",x"9E"),
		(x"01",x"05",x"05",x"06",x"00",x"00",x"00",x"07",x"07",x"03",x"03",x"07",x"00",x"07",x"04",x"00",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"00",x"09",x"00",x"0D",x"01",x"08",x"09"),
		(x"04",x"01",x"04",x"00",x"0C",x"0E",x"04",x"05",x"03",x"01",x"03",x"00",x"16",x"04",x"04",x"0E",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"0A",x"00",x"05",x"07",x"00",x"03",x"00"),
		(x"01",x"00",x"07",x"A1",x"A4",x"A4",x"1E",x"1A",x"A3",x"A2",x"A7",x"A1",x"A2",x"1D",x"A6",x"A0",x"1C",x"1C",x"1C",x"1C",x"1C",x"1C",x"1C",x"1C",x"9A",x"1B",x"A6",x"A9",x"98",x"0F",x"08"),
		(x"01",x"00",x"07",x"A1",x"A4",x"A4",x"1E",x"1A",x"A3",x"A2",x"A7",x"A1",x"A2",x"1D",x"A6",x"A0",x"1C",x"1C",x"1C",x"1C",x"1C",x"1C",x"1C",x"1C",x"21",x"AA",x"19",x"A8",x"9E",x"0B",x"00"),
		(x"01",x"00",x"07",x"A1",x"A4",x"A4",x"1E",x"1A",x"A3",x"A2",x"A7",x"A1",x"A2",x"1D",x"A6",x"A0",x"1C",x"1C",x"1C",x"1C",x"1C",x"1C",x"1C",x"1C",x"9A",x"20",x"A0",x"A8",x"99",x"0B",x"00"),
		(x"01",x"00",x"07",x"A1",x"A4",x"A4",x"1E",x"1A",x"A3",x"A2",x"A7",x"A1",x"A2",x"1D",x"A6",x"A0",x"1C",x"1C",x"1C",x"1C",x"1C",x"1C",x"1C",x"1C",x"18",x"A9",x"14",x"9E",x"A1",x"0A",x"00"),
		(x"01",x"00",x"07",x"A1",x"A4",x"A4",x"1E",x"1A",x"A3",x"A2",x"A7",x"A1",x"A2",x"1D",x"A6",x"A0",x"1C",x"1C",x"1C",x"1C",x"1C",x"1C",x"1C",x"1C",x"A0",x"21",x"A6",x"AC",x"A3",x"03",x"09"),
		(x"01",x"00",x"07",x"A1",x"A4",x"A4",x"1E",x"1A",x"A3",x"A2",x"A7",x"A1",x"A2",x"1D",x"A6",x"A0",x"1C",x"1C",x"1C",x"1C",x"1C",x"1C",x"1C",x"1C",x"1E",x"AA",x"19",x"A1",x"AA",x"03",x"06"),
		(x"01",x"00",x"07",x"A1",x"A4",x"A4",x"1E",x"1A",x"A3",x"A2",x"A7",x"A1",x"A2",x"1D",x"A6",x"A0",x"1C",x"1C",x"1C",x"1C",x"1C",x"1C",x"1C",x"1C",x"98",x"1F",x"A1",x"A0",x"A5",x"02",x"07"),
		(x"01",x"00",x"07",x"A1",x"A4",x"A4",x"1E",x"1A",x"A3",x"A2",x"A7",x"A1",x"A2",x"1D",x"A6",x"A0",x"1C",x"1C",x"1C",x"1C",x"1C",x"1C",x"1C",x"1C",x"1E",x"AF",x"15",x"9F",x"AB",x"00",x"00"),
		(x"01",x"00",x"07",x"A1",x"A4",x"A4",x"1E",x"1A",x"A3",x"A2",x"A7",x"A1",x"A2",x"1D",x"A6",x"A0",x"1C",x"1C",x"1C",x"1C",x"1C",x"1C",x"1C",x"1C",x"9A",x"1B",x"A6",x"A9",x"98",x"0F",x"08"),
		(x"01",x"00",x"07",x"A1",x"A4",x"A4",x"1E",x"1A",x"A3",x"A2",x"A7",x"A1",x"A2",x"1D",x"A6",x"A0",x"1C",x"1C",x"1C",x"1C",x"1C",x"1C",x"1C",x"1C",x"21",x"AA",x"19",x"A8",x"9E",x"0B",x"00"),
		(x"01",x"00",x"07",x"A1",x"A4",x"A4",x"1E",x"1A",x"A3",x"A2",x"A7",x"A1",x"A2",x"1D",x"A6",x"A0",x"1C",x"1C",x"1C",x"1C",x"1C",x"1C",x"1C",x"1C",x"9A",x"20",x"A0",x"A8",x"99",x"0B",x"00"),
		(x"01",x"00",x"07",x"A1",x"A4",x"A4",x"1E",x"1A",x"A3",x"A2",x"A7",x"A1",x"A2",x"1D",x"A6",x"A0",x"1C",x"1C",x"1C",x"1C",x"1C",x"1C",x"1C",x"1C",x"18",x"A9",x"14",x"9E",x"A1",x"0A",x"00"),
		(x"01",x"00",x"07",x"A1",x"A4",x"A4",x"1E",x"1A",x"A3",x"A2",x"A7",x"A1",x"A2",x"1D",x"A6",x"A0",x"1C",x"1C",x"1C",x"1C",x"1C",x"1C",x"1C",x"1C",x"A0",x"21",x"A6",x"AC",x"A3",x"03",x"09"),
		(x"01",x"00",x"07",x"A1",x"A4",x"A4",x"1E",x"1A",x"A3",x"A2",x"A7",x"A1",x"A2",x"1D",x"A6",x"A0",x"1C",x"1C",x"1C",x"1C",x"1C",x"1C",x"1C",x"1C",x"1E",x"AA",x"19",x"A1",x"AA",x"03",x"06"),
		(x"01",x"00",x"07",x"A1",x"A4",x"A4",x"1E",x"1A",x"A3",x"A2",x"A7",x"A1",x"A2",x"1D",x"A6",x"A0",x"1C",x"1C",x"1C",x"1C",x"1C",x"1C",x"1C",x"1C",x"98",x"1F",x"A1",x"A0",x"A5",x"02",x"07")
	
	);
	
	constant pipe_G : ROM :=
	(
	
		(x"09",x"00",x"05",x"04",x"09",x"00",x"0A",x"01",x"0C",x"08",x"06",x"09",x"04",x"05",x"03",x"00",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"08",x"00",x"05",x"09",x"00",x"08",x"00"),
		(x"00",x"B9",x"C2",x"B5",x"C0",x"C4",x"B6",x"C3",x"B5",x"B4",x"BA",x"BE",x"B2",x"BF",x"C3",x"BD",x"BC",x"BC",x"BC",x"BC",x"BC",x"BC",x"BC",x"BC",x"BD",x"BE",x"BA",x"BC",x"C4",x"BF",x"B3"),
		(x"14",x"79",x"7D",x"87",x"88",x"76",x"C3",x"B3",x"BF",x"B9",x"BD",x"BB",x"86",x"80",x"85",x"81",x"83",x"83",x"83",x"83",x"83",x"83",x"83",x"83",x"81",x"93",x"78",x"82",x"7B",x"88",x"8C"),
		(x"00",x"C5",x"B6",x"C1",x"83",x"8A",x"C1",x"B8",x"BE",x"BF",x"BC",x"B5",x"8F",x"BD",x"BB",x"87",x"85",x"85",x"85",x"85",x"85",x"85",x"85",x"85",x"7E",x"BF",x"82",x"BC",x"86",x"BD",x"BB"),
		(x"00",x"BB",x"BA",x"B6",x"84",x"7A",x"BA",x"BB",x"C0",x"BA",x"BA",x"BE",x"8B",x"B9",x"B8",x"89",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"7F",x"88",x"7A",x"B9",x"87",x"B7",x"C3",x"B9"),
		(x"07",x"C6",x"C1",x"BA",x"84",x"8D",x"BE",x"BD",x"B3",x"BD",x"BD",x"B6",x"7C",x"BF",x"BD",x"7F",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"87",x"85",x"C5",x"82",x"C0",x"76",x"BF",x"B3"),
		(x"00",x"B9",x"BF",x"C0",x"77",x"7F",x"B7",x"C6",x"C0",x"BF",x"BB",x"C3",x"86",x"BA",x"B7",x"8A",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"7D",x"88",x"BA",x"85",x"C6",x"B5",x"C8"),
		(x"0B",x"B2",x"BD",x"C3",x"83",x"8A",x"BE",x"B2",x"BB",x"BD",x"B7",x"BC",x"84",x"C0",x"BA",x"85",x"83",x"83",x"83",x"83",x"83",x"83",x"83",x"83",x"87",x"B8",x"84",x"C0",x"7E",x"BF",x"C2"),
		(x"0B",x"C4",x"B3",x"BD",x"7F",x"8D",x"BF",x"BA",x"C0",x"B9",x"BD",x"BD",x"7E",x"C0",x"C5",x"7B",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"85",x"7A",x"C3",x"87",x"BC",x"BD",x"B9"),
		(x"04",x"B2",x"BC",x"BD",x"83",x"8E",x"B1",x"C0",x"B9",x"BC",x"BA",x"B5",x"87",x"BD",x"BC",x"83",x"83",x"83",x"83",x"83",x"83",x"83",x"83",x"83",x"83",x"BB",x"7F",x"B4",x"80",x"B9",x"B9"),
		(x"02",x"C4",x"BA",x"BE",x"84",x"7E",x"BC",x"BA",x"C1",x"B8",x"C5",x"BE",x"7C",x"BB",x"C8",x"78",x"85",x"85",x"85",x"85",x"85",x"85",x"85",x"85",x"8A",x"83",x"BA",x"89",x"BC",x"BF",x"B1"),
		(x"06",x"B7",x"B6",x"BF",x"87",x"81",x"B6",x"C2",x"BE",x"B6",x"B8",x"BE",x"87",x"BB",x"BC",x"87",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"81",x"C1",x"7F",x"BF",x"8C",x"AE",x"C5"),
		(x"03",x"BE",x"BE",x"BE",x"83",x"89",x"BD",x"B4",x"BB",x"BF",x"BB",x"BA",x"83",x"C0",x"BC",x"82",x"83",x"83",x"83",x"83",x"83",x"83",x"83",x"83",x"83",x"7A",x"C1",x"7C",x"BE",x"BB",x"BE"),
		(x"0C",x"B8",x"BC",x"BA",x"79",x"7B",x"C2",x"BD",x"BB",x"BB",x"BC",x"BB",x"84",x"BD",x"BE",x"84",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"82",x"7F",x"C4",x"89",x"AF",x"87",x"C0",x"B7"),
		(x"02",x"07",x"00",x"09",x"0A",x"0E",x"05",x"00",x"07",x"06",x"01",x"0A",x"06",x"06",x"00",x"09",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"09",x"03",x"01",x"0A",x"02",x"02",x"09"),
		(x"00",x"00",x"09",x"05",x"01",x"00",x"05",x"04",x"02",x"06",x"08",x"01",x"04",x"01",x"03",x"04",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"03",x"02",x"08",x"05",x"00",x"0B",x"01",x"05"),
		(x"00",x"02",x"04",x"BB",x"BE",x"BB",x"84",x"84",x"BD",x"BC",x"BB",x"BC",x"BC",x"85",x"B8",x"BE",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"BD",x"86",x"BB",x"BC",x"BF",x"05",x"00"),
		(x"00",x"02",x"04",x"BB",x"BE",x"BB",x"84",x"84",x"BD",x"BC",x"BB",x"BC",x"BC",x"85",x"B8",x"BE",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"86",x"BA",x"81",x"BC",x"BD",x"01",x"08"),
		(x"00",x"02",x"04",x"BB",x"BE",x"BB",x"84",x"84",x"BD",x"BC",x"BB",x"BC",x"BC",x"85",x"B8",x"BE",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"BD",x"7C",x"C8",x"B3",x"BE",x"07",x"00"),
		(x"00",x"02",x"04",x"BB",x"BE",x"BB",x"84",x"84",x"BD",x"BC",x"BB",x"BC",x"BC",x"85",x"B8",x"BE",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"8A",x"BA",x"80",x"C3",x"B9",x"08",x"01"),
		(x"00",x"02",x"04",x"BB",x"BE",x"BB",x"84",x"84",x"BD",x"BC",x"BB",x"BC",x"BC",x"85",x"B8",x"BE",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"BA",x"81",x"C1",x"B8",x"BD",x"02",x"04"),
		(x"00",x"02",x"04",x"BB",x"BE",x"BB",x"84",x"84",x"BD",x"BC",x"BB",x"BC",x"BC",x"85",x"B8",x"BE",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"87",x"BF",x"78",x"C7",x"B8",x"04",x"02"),
		(x"00",x"02",x"04",x"BB",x"BE",x"BB",x"84",x"84",x"BD",x"BC",x"BB",x"BC",x"BC",x"85",x"B8",x"BE",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"BF",x"82",x"BF",x"BE",x"B9",x"08",x"00"),
		(x"00",x"02",x"04",x"BB",x"BE",x"BB",x"84",x"84",x"BD",x"BC",x"BB",x"BC",x"BC",x"85",x"B8",x"BE",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"88",x"B5",x"85",x"BE",x"B7",x"04",x"07"),
		(x"00",x"02",x"04",x"BB",x"BE",x"BB",x"84",x"84",x"BD",x"BC",x"BB",x"BC",x"BC",x"85",x"B8",x"BE",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"BD",x"86",x"BB",x"BC",x"BF",x"05",x"00"),
		(x"00",x"02",x"04",x"BB",x"BE",x"BB",x"84",x"84",x"BD",x"BC",x"BB",x"BC",x"BC",x"85",x"B8",x"BE",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"86",x"BA",x"81",x"BC",x"BD",x"01",x"08"),
		(x"00",x"02",x"04",x"BB",x"BE",x"BB",x"84",x"84",x"BD",x"BC",x"BB",x"BC",x"BC",x"85",x"B8",x"BE",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"BD",x"7C",x"C8",x"B3",x"BE",x"07",x"00"),
		(x"00",x"02",x"04",x"BB",x"BE",x"BB",x"84",x"84",x"BD",x"BC",x"BB",x"BC",x"BC",x"85",x"B8",x"BE",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"8A",x"BA",x"80",x"C3",x"B9",x"08",x"01"),
		(x"00",x"02",x"04",x"BB",x"BE",x"BB",x"84",x"84",x"BD",x"BC",x"BB",x"BC",x"BC",x"85",x"B8",x"BE",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"BA",x"81",x"C1",x"B8",x"BD",x"02",x"04"),
		(x"00",x"02",x"04",x"BB",x"BE",x"BB",x"84",x"84",x"BD",x"BC",x"BB",x"BC",x"BC",x"85",x"B8",x"BE",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"87",x"BF",x"78",x"C7",x"B8",x"04",x"02"),
		(x"00",x"02",x"04",x"BB",x"BE",x"BB",x"84",x"84",x"BD",x"BC",x"BB",x"BC",x"BC",x"85",x"B8",x"BE",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"BF",x"82",x"BF",x"BE",x"B9",x"08",x"00")
	
	);
	
	constant pipe_B : ROM :=
	(
	
		(x"0B",x"02",x"04",x"00",x"04",x"09",x"0D",x"0A",x"05",x"01",x"04",x"0F",x"00",x"01",x"07",x"02",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"00",x"0E",x"01",x"03",x"0B",x"07",x"00"),
		(x"05",x"07",x"00",x"16",x"00",x"00",x"00",x"00",x"00",x"00",x"02",x"00",x"00",x"05",x"09",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"05",x"01",x"00",x"00",x"00",x"00",x"05"),
		(x"02",x"19",x"18",x"06",x"1B",x"10",x"15",x"07",x"12",x"00",x"00",x"00",x"1E",x"1B",x"15",x"0B",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"0F",x"13",x"17",x"1E",x"17",x"1B",x"1B"),
		(x"04",x"04",x"00",x"0E",x"16",x"1A",x"00",x"00",x"00",x"00",x"0A",x"02",x"14",x"00",x"0B",x"1A",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"14",x"0C",x"11",x"03",x"20",x"00",x"04"),
		(x"0A",x"00",x"00",x"14",x"14",x"0B",x"03",x"04",x"0A",x"00",x"04",x"04",x"16",x"00",x"00",x"10",x"1B",x"1B",x"1B",x"1B",x"1B",x"1B",x"1B",x"1B",x"07",x"17",x"04",x"14",x"00",x"00",x"0C"),
		(x"09",x"0F",x"00",x"00",x"26",x"14",x"00",x"00",x"00",x"08",x"07",x"00",x"0E",x"0D",x"0B",x"09",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"09",x"04",x"1A",x"00",x"2B",x"00",x"01"),
		(x"00",x"0A",x"00",x"00",x"23",x"1B",x"00",x"00",x"00",x"00",x"00",x"00",x"0B",x"0A",x"07",x"13",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"16",x"0F",x"0D",x"00",x"03",x"11",x"07",x"00"),
		(x"00",x"07",x"00",x"00",x"1A",x"01",x"0B",x"0A",x"0B",x"09",x"00",x"0D",x"0E",x"07",x"00",x"0F",x"15",x"15",x"15",x"15",x"15",x"15",x"15",x"15",x"1E",x"08",x"24",x"00",x"17",x"02",x"0C"),
		(x"00",x"14",x"02",x"05",x"0F",x"00",x"06",x"00",x"00",x"00",x"00",x"04",x"17",x"00",x"00",x"21",x"15",x"15",x"15",x"15",x"15",x"15",x"15",x"15",x"12",x"15",x"04",x"1B",x"00",x"00",x"10"),
		(x"00",x"01",x"07",x"00",x"17",x"1C",x"05",x"00",x"00",x"09",x"00",x"00",x"1E",x"00",x"00",x"22",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"1B",x"01",x"11",x"00",x"10",x"08",x"00"),
		(x"00",x"0C",x"07",x"00",x"0E",x"17",x"0D",x"00",x"04",x"00",x"0F",x"04",x"0F",x"00",x"09",x"0C",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"1F",x"17",x"00",x"15",x"09",x"03",x"01"),
		(x"0A",x"00",x"00",x"00",x"14",x"22",x"00",x"00",x"01",x"00",x"00",x"00",x"1B",x"00",x"00",x"19",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"13",x"04",x"06",x"1F",x"00",x"19",x"0A",x"01"),
		(x"08",x"07",x"00",x"12",x"14",x"20",x"00",x"00",x"00",x"06",x"00",x"00",x"1B",x"07",x"00",x"18",x"15",x"15",x"15",x"15",x"15",x"15",x"15",x"15",x"1E",x"08",x"00",x"21",x"08",x"04",x"00"),
		(x"00",x"00",x"00",x"06",x"09",x"15",x"06",x"00",x"04",x"04",x"00",x"04",x"08",x"09",x"04",x"08",x"15",x"15",x"15",x"15",x"15",x"15",x"15",x"15",x"16",x"00",x"2B",x"00",x"15",x"00",x"04"),
		(x"17",x"02",x"0A",x"12",x"05",x"05",x"00",x"11",x"00",x"00",x"00",x"03",x"0E",x"01",x"00",x"12",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"11",x"07",x"0E",x"01",x"00",x"0C",x"09"),
		(x"00",x"00",x"05",x"00",x"00",x"0D",x"0A",x"09",x"07",x"0A",x"0E",x"07",x"00",x"08",x"0B",x"00",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"05",x"00",x"03",x"00",x"0C",x"02",x"0F",x"00"),
		(x"02",x"02",x"00",x"04",x"03",x"00",x"14",x"16",x"00",x"05",x"01",x"00",x"01",x"16",x"00",x"00",x"15",x"15",x"15",x"15",x"15",x"15",x"15",x"15",x"01",x"26",x"00",x"0A",x"00",x"06",x"00"),
		(x"02",x"02",x"00",x"04",x"03",x"00",x"14",x"16",x"00",x"05",x"01",x"00",x"01",x"16",x"00",x"00",x"15",x"15",x"15",x"15",x"15",x"15",x"15",x"15",x"04",x"02",x"0E",x"00",x"00",x"02",x"0A"),
		(x"02",x"02",x"00",x"04",x"03",x"00",x"14",x"16",x"00",x"05",x"01",x"00",x"01",x"16",x"00",x"00",x"15",x"15",x"15",x"15",x"15",x"15",x"15",x"15",x"00",x"19",x"07",x"00",x"00",x"08",x"05"),
		(x"02",x"02",x"00",x"04",x"03",x"00",x"14",x"16",x"00",x"05",x"01",x"00",x"01",x"16",x"00",x"00",x"15",x"15",x"15",x"15",x"15",x"15",x"15",x"15",x"18",x"00",x"1D",x"03",x"01",x"0B",x"02"),
		(x"02",x"02",x"00",x"04",x"03",x"00",x"14",x"16",x"00",x"05",x"01",x"00",x"01",x"16",x"00",x"00",x"15",x"15",x"15",x"15",x"15",x"15",x"15",x"15",x"00",x"1F",x"00",x"00",x"00",x"00",x"08"),
		(x"02",x"02",x"00",x"04",x"03",x"00",x"14",x"16",x"00",x"05",x"01",x"00",x"01",x"16",x"00",x"00",x"15",x"15",x"15",x"15",x"15",x"15",x"15",x"15",x"10",x"00",x"10",x"02",x"00",x"00",x"01"),
		(x"02",x"02",x"00",x"04",x"03",x"00",x"14",x"16",x"00",x"05",x"01",x"00",x"01",x"16",x"00",x"00",x"15",x"15",x"15",x"15",x"15",x"15",x"15",x"15",x"0A",x"16",x"09",x"04",x"00",x"04",x"00"),
		(x"02",x"02",x"00",x"04",x"03",x"00",x"14",x"16",x"00",x"05",x"01",x"00",x"01",x"16",x"00",x"00",x"15",x"15",x"15",x"15",x"15",x"15",x"15",x"15",x"0E",x"00",x"23",x"00",x"00",x"02",x"18"),
		(x"02",x"02",x"00",x"04",x"03",x"00",x"14",x"16",x"00",x"05",x"01",x"00",x"01",x"16",x"00",x"00",x"15",x"15",x"15",x"15",x"15",x"15",x"15",x"15",x"01",x"26",x"00",x"0A",x"00",x"06",x"00"),
		(x"02",x"02",x"00",x"04",x"03",x"00",x"14",x"16",x"00",x"05",x"01",x"00",x"01",x"16",x"00",x"00",x"15",x"15",x"15",x"15",x"15",x"15",x"15",x"15",x"04",x"02",x"0E",x"00",x"00",x"02",x"0A"),
		(x"02",x"02",x"00",x"04",x"03",x"00",x"14",x"16",x"00",x"05",x"01",x"00",x"01",x"16",x"00",x"00",x"15",x"15",x"15",x"15",x"15",x"15",x"15",x"15",x"00",x"19",x"07",x"00",x"00",x"08",x"05"),
		(x"02",x"02",x"00",x"04",x"03",x"00",x"14",x"16",x"00",x"05",x"01",x"00",x"01",x"16",x"00",x"00",x"15",x"15",x"15",x"15",x"15",x"15",x"15",x"15",x"18",x"00",x"1D",x"03",x"01",x"0B",x"02"),
		(x"02",x"02",x"00",x"04",x"03",x"00",x"14",x"16",x"00",x"05",x"01",x"00",x"01",x"16",x"00",x"00",x"15",x"15",x"15",x"15",x"15",x"15",x"15",x"15",x"00",x"1F",x"00",x"00",x"00",x"00",x"08"),
		(x"02",x"02",x"00",x"04",x"03",x"00",x"14",x"16",x"00",x"05",x"01",x"00",x"01",x"16",x"00",x"00",x"15",x"15",x"15",x"15",x"15",x"15",x"15",x"15",x"10",x"00",x"10",x"02",x"00",x"00",x"01"),
		(x"02",x"02",x"00",x"04",x"03",x"00",x"14",x"16",x"00",x"05",x"01",x"00",x"01",x"16",x"00",x"00",x"15",x"15",x"15",x"15",x"15",x"15",x"15",x"15",x"0A",x"16",x"09",x"04",x"00",x"04",x"00")
	
	);
	
begin

	dat_R <= pipe_R( dir_y )( dir_x );
	dat_G <= pipe_G( dir_y )( dir_x );
	dat_B <= pipe_B( dir_y )( dir_x );

end comp;