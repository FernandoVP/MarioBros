library ieee;

use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity bg4_ROM is

	Port(
	
		dir_y : in integer;
		dir_x : in integer;
		
		dat_R : out std_logic_vector( 7 downto 0 );
		dat_G : out std_logic_vector( 7 downto 0 );
		dat_B : out std_logic_vector( 7 downto 0 )
		
	);

end bg4_ROM;

architecture comp of bg4_ROM is

	type arreglo is array( 0 to 119 ) of std_logic_vector( 0 to 7 );

	type ROM is array( 0 to 76 ) of arreglo;

	constant bg_R : ROM :=
	(
	
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"EF",x"EF",x"EF",x"EF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"EF",x"EF",x"EF",x"EF",x"EF",x"EF",x"EF",x"EF",x"EF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"EF",x"EF",x"EF",x"EF",x"EF",x"EF",x"EF",x"EF",x"EF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"EF",x"EF",x"EF",x"EF",x"EF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"E9",x"E9",x"E9",x"F0",x"01",x"00",x"00",x"00",x"01",x"00",x"00",x"EF",x"E8",x"E9",x"E7",x"E8",x"E9",x"E8",x"E9",x"F0",x"01",x"00",x"00",x"00",x"01",x"00",x"00",x"EF",x"E8",x"E9",x"E7",x"E8",x"E9",x"E8",x"E9",x"F0",x"01",x"00",x"00",x"00",x"01",x"00",x"00",x"EF",x"E8",x"E8",x"E8",x"E8",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E9",x"E8",x"E8",x"F7",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"F0",x"E8",x"E8",x"E8",x"E8",x"E9",x"E8",x"E8",x"F7",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"F0",x"E8",x"E8",x"E8",x"E8",x"E9",x"E8",x"E8",x"F7",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"F0",x"E8",x"E8",x"E8",x"E8",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E8",x"E7",x"E8",x"EF",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"EF",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"EE",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"EF",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"EE",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"EF",x"E8",x"E8",x"E8",x"E8",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E8",x"E8",x"E8",x"F7",x"00",x"01",x"00",x"00",x"01",x"00",x"00",x"EF",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"F7",x"00",x"01",x"00",x"00",x"01",x"00",x"00",x"EF",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"F7",x"00",x"01",x"00",x"00",x"01",x"00",x"00",x"EF",x"E8",x"E8",x"E8",x"E8",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E8",x"E8",x"E8",x"EF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"EF",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"EF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"EF",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"EF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"EF",x"E8",x"E8",x"E8",x"E8",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E8",x"E8",x"E9",x"F7",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"EF",x"E8",x"E9",x"E8",x"E7",x"E9",x"E9",x"E9",x"F7",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"EF",x"E8",x"E9",x"E8",x"E7",x"E9",x"E9",x"E9",x"F7",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"EF",x"E8",x"E8",x"E8",x"E8",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"F0",x"EF",x"EF",x"EF",x"EF",x"EF",x"EF",x"EF",x"EF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"EF",x"EF",x"EF",x"EF",x"EF",x"EF",x"EF",x"EF",x"EF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"EF",x"EF",x"EF",x"EF",x"EF",x"EF",x"EF",x"EF",x"EF",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E8",x"E8",x"E9",x"E7",x"E7",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"E8",x"E9",x"E8",x"E8",x"E7",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"E8",x"E9",x"E8",x"E8",x"E7",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E8",x"E9",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E9",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"E7",x"00",x"E8",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"E7",x"00",x"E8",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"E8",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"01",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"01",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"E9",x"00",x"E8",x"E8",x"E8",x"E8",x"E9",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"E9",x"00",x"E8",x"E8",x"E8",x"E8",x"E9",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"E9",x"00",x"E6",x"E8",x"E7",x"E8",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E7",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"E9",x"00",x"E8",x"E8",x"E8",x"E9",x"E7",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"E9",x"00",x"E8",x"E8",x"E8",x"E9",x"E7",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"E9",x"00",x"E8",x"E8",x"E8",x"E8",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E8",x"E8",x"E8",x"E7",x"E8",x"E8",x"E8",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"E8",x"E8",x"E8",x"E7",x"E8",x"E8",x"E8",x"00",x"E9",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"E8",x"E8",x"E8",x"E7",x"E8",x"E8",x"E8",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"E8",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"E8",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"00",x"E7",x"E8",x"E8",x"E8",x"E7",x"E8",x"E8",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"E8",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"E8",x"E8",x"E8",x"00",x"E6",x"E8",x"E7",x"E8",x"00",x"00",x"01",x"00",x"00",x"01",x"00",x"00",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"E8",x"00",x"E6",x"E8",x"E7",x"E8",x"00",x"00",x"01",x"00",x"00",x"01",x"00",x"00",x"E8",x"E8",x"E8",x"00",x"E6",x"E8",x"E7",x"E8",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E9",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E9",x"E8",x"E8",x"00",x"E9",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E9",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E9",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E8",x"E8",x"E8",x"E7",x"E8",x"E8",x"E8",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"E8",x"E8",x"E8",x"E7",x"E8",x"E8",x"E8",x"00",x"E9",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"E8",x"E8",x"E8",x"E7",x"E8",x"E8",x"E8",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"E8",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"E8",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"00",x"E7",x"E8",x"E8",x"E8",x"E7",x"E8",x"E8",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"E8",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"E8",x"E8",x"E8",x"00",x"E6",x"E8",x"E7",x"E8",x"00",x"00",x"01",x"00",x"00",x"01",x"00",x"00",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"E8",x"00",x"E6",x"E8",x"E7",x"E8",x"00",x"00",x"01",x"00",x"00",x"01",x"00",x"00",x"E8",x"E8",x"E8",x"00",x"E6",x"E8",x"E7",x"E8",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E9",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E9",x"E8",x"E8",x"00",x"E9",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E9",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E9",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"EF",x"EF",x"EF",x"EF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"EF",x"EF",x"EF",x"EF",x"EF",x"EF",x"EF",x"F0",x"EF",x"E8",x"E8",x"E9",x"00",x"E8",x"E8",x"E8",x"EF",x"EF",x"EF",x"EF",x"EF",x"EF",x"EF",x"EF",x"EF",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"F7",x"EF",x"EF",x"F7",x"EF",x"EF",x"EF",x"EF",x"EF",x"E8",x"E9",x"E8",x"00",x"E8",x"E8",x"E7",x"F7",x"EF",x"EF",x"F7",x"EF",x"EF",x"EF",x"EF",x"EE",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"EF",x"EF",x"EF",x"EF",x"EF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"E9",x"E9",x"E9",x"F0",x"01",x"00",x"00",x"00",x"01",x"00",x"00",x"EF",x"E8",x"E9",x"E8",x"E8",x"E9",x"E8",x"E9",x"F7",x"E7",x"E8",x"E8",x"00",x"E8",x"E7",x"E8",x"F7",x"E8",x"E9",x"E7",x"E8",x"E9",x"E8",x"E9",x"F0",x"E7",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"F7",x"E8",x"E9",x"E8",x"E8",x"E9",x"E8",x"E9",x"EF",x"E7",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"EF",x"E8",x"E9",x"E8",x"E8",x"E9",x"E8",x"E9",x"EF",x"01",x"00",x"00",x"00",x"01",x"00",x"00",x"EF",x"E8",x"E8",x"E8",x"E8",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E9",x"E8",x"E8",x"F7",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"F0",x"E8",x"E8",x"E8",x"E8",x"E9",x"E8",x"E8",x"EF",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"F7",x"E8",x"E8",x"E8",x"E8",x"E9",x"E8",x"E8",x"F7",x"E8",x"E9",x"E8",x"00",x"E8",x"E8",x"E8",x"EF",x"E8",x"E9",x"E8",x"E8",x"E8",x"E8",x"E8",x"F7",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"F7",x"E8",x"E8",x"E8",x"E8",x"E9",x"E8",x"E8",x"EF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"F0",x"E8",x"E8",x"E8",x"E8",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E8",x"E7",x"E8",x"EF",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"EF",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"F7",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"F0",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"EE",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"F9",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"EF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"F0",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"F8",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"EF",x"E8",x"E8",x"E8",x"E8",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E8",x"E8",x"E8",x"F7",x"00",x"01",x"00",x"00",x"01",x"00",x"00",x"EF",x"E9",x"E8",x"E8",x"E8",x"E9",x"E8",x"E8",x"F7",x"E8",x"E8",x"E8",x"E8",x"E9",x"E8",x"E8",x"EF",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"F7",x"E8",x"E8",x"E8",x"E8",x"E9",x"E8",x"E8",x"EF",x"E8",x"E7",x"E8",x"E7",x"E8",x"E8",x"E8",x"F7",x"E8",x"E8",x"E9",x"E8",x"E9",x"E8",x"E8",x"EF",x"E9",x"E8",x"E8",x"E8",x"E8",x"E9",x"E7",x"EF",x"00",x"01",x"00",x"00",x"01",x"00",x"00",x"EF",x"E8",x"E8",x"E8",x"E8",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E8",x"E8",x"E8",x"EF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"EF",x"E8",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"EF",x"E8",x"E9",x"E8",x"E9",x"E8",x"E8",x"E8",x"F7",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"EF",x"E8",x"E9",x"E8",x"EA",x"E9",x"E8",x"E9",x"F7",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"EF",x"E8",x"E9",x"E9",x"E8",x"E8",x"E8",x"E8",x"F8",x"E8",x"E8",x"E7",x"E8",x"E8",x"E9",x"E8",x"F7",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"EF",x"E8",x"E8",x"E8",x"E8",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E8",x"E8",x"E9",x"F7",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"EF",x"E8",x"E9",x"E8",x"E7",x"E8",x"E8",x"E9",x"F7",x"E8",x"E8",x"E7",x"E8",x"E8",x"E9",x"E8",x"EF",x"E8",x"E9",x"E8",x"E7",x"E9",x"E9",x"E9",x"F7",x"E8",x"E8",x"E7",x"E8",x"E9",x"E8",x"E8",x"EF",x"E8",x"E9",x"E8",x"E7",x"E7",x"E8",x"E9",x"F7",x"E8",x"E8",x"E7",x"E8",x"E8",x"E8",x"E8",x"EF",x"E8",x"E9",x"E8",x"E7",x"E8",x"E8",x"E9",x"EF",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"EF",x"E8",x"E8",x"E8",x"E8",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"F0",x"EF",x"EF",x"EF",x"EF",x"EF",x"EF",x"EF",x"EF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"EF",x"F6",x"EF",x"F7",x"EF",x"F7",x"EF",x"F7",x"EF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"EF",x"F6",x"EF",x"F7",x"EF",x"F7",x"EF",x"F7",x"EF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"EF",x"F6",x"EF",x"F7",x"EF",x"F7",x"EF",x"F7",x"EF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"F7",x"EF",x"EF",x"EF",x"EF",x"EF",x"EF",x"EF",x"EF",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E8",x"E8",x"E9",x"E7",x"E7",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"E8",x"E9",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"E8",x"E9",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"E8",x"E9",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E8",x"E9",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E8",x"E9",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"00",x"E9",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"00",x"E9",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"00",x"E9",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E9",x"E8",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E9",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"E7",x"00",x"E8",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"00",x"E8",x"E8",x"E8",x"E9",x"E8",x"E8",x"E7",x"00",x"E8",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"00",x"E8",x"E8",x"E8",x"E9",x"E8",x"E8",x"E7",x"00",x"E8",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"00",x"E8",x"E8",x"E8",x"E9",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E7",x"E8",x"E8",x"E7",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"E8",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"01",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"01",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"01",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"01",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"E9",x"00",x"E8",x"E8",x"E8",x"E8",x"E9",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E9",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E9",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E9",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"E9",x"00",x"E6",x"E8",x"E7",x"E8",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E7",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"E9",x"00",x"E8",x"E8",x"E8",x"E9",x"E7",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"E9",x"00",x"E8",x"E8",x"E8",x"E9",x"E7",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"E9",x"00",x"E8",x"E8",x"E8",x"E9",x"E7",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"E9",x"00",x"E8",x"E8",x"E8",x"E9",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"E9",x"00",x"E8",x"E8",x"E8",x"E8",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E8",x"E7",x"E8",x"E8",x"E7",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E9",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E9",x"00",x"00",x"00",x"00",x"00",x"00",x"E9",x"E8",x"E8",x"E8",x"00",x"E7",x"E9",x"E9",x"E8",x"E7",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E8",x"E8",x"E8",x"E7",x"E8",x"E8",x"E8",x"00",x"E9",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"E9",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"E9",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"E8",x"E7",x"E8",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E8",x"E8",x"00",x"E8",x"E7",x"E7",x"E8",x"E8",x"E8",x"E8",x"00",x"E9",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"E9",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"E9",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"BD",x"BD",x"BD",x"BD",x"00",x"00",x"01",x"00",x"00",x"01",x"E8",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"00",x"E7",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"00",x"E7",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"00",x"E7",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"00",x"E8",x"E8",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E8",x"01",x"E7",x"E8",x"E8",x"E9",x"E8",x"E7",x"E8",x"00",x"E7",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"00",x"E7",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"00",x"E7",x"E8",x"E8",x"E8",x"E7",x"E8",x"E8",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"BD",x"BD",x"FE",x"FE",x"FE",x"FE",x"BD",x"BD",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"BD",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"BD",x"01",x"00",x"00",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"E8",x"00",x"E7",x"E7",x"E8",x"E8",x"E8",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E8",x"E8",x"E9",x"E9",x"00",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"E8",x"00",x"E6",x"E8",x"E7",x"E8",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"BE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"BD",x"00",x"00",x"E9",x"E8",x"E8",x"00",x"E9",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"E9",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"E9",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E8",x"E8",x"E8",x"E9",x"00",x"E9",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"E9",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"E9",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"BD",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FF",x"BC",x"01",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E9",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E9",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E9",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E7",x"E9",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"E7",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E9",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E9",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E9",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"01",x"00",x"00",x"00",x"BD",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"BD",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"BE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FF",x"FE",x"BD",x"00",x"E8",x"E8",x"E8",x"E9",x"E7",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"BD",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"BD",x"00",x"E8",x"E8",x"E8",x"E7",x"E8",x"E8",x"E8",x"00",x"E9",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"E9",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"E9",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E8",x"E8",x"E8",x"E7",x"E8",x"E8",x"E8",x"00",x"E9",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"E9",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"E9",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"BD",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FF",x"FE",x"BD",x"00",x"E8",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"00",x"E7",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"00",x"E7",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"00",x"E7",x"E8",x"E8",x"E8",x"E7",x"E8",x"E8",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"E8",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"00",x"E7",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"00",x"E7",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"00",x"E7",x"E8",x"E8",x"E8",x"E7",x"E8",x"E8",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"BD",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"BD",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"01",x"00",x"00",x"BE",x"BD",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"BD",x"BE",x"00",x"00",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"E8",x"00",x"E6",x"E8",x"E7",x"E8",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"E8",x"00",x"E6",x"E8",x"E7",x"E8",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"BD",x"BD",x"BD",x"FE",x"FE",x"FE",x"FE",x"BD",x"BD",x"BD",x"00",x"00",x"00",x"E9",x"E8",x"E8",x"00",x"E9",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"E9",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"E9",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E9",x"E8",x"E8",x"00",x"E9",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"E9",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"E9",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"BD",x"BD",x"BD",x"BD",x"BD",x"BD",x"BD",x"BD",x"00",x"00",x"00",x"01",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E9",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E9",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E9",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E9",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E9",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E9",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"BD",x"BE",x"BC",x"BD",x"BC",x"C7",x"BE",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"EF",x"F7",x"EF",x"F0",x"F7",x"EF",x"00",x"00",x"00",x"00",x"00",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"01",x"00",x"00",x"00",x"EF",x"E8",x"ED",x"EF",x"EF",x"E8",x"E8",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"EF",x"EF",x"EF",x"F0",x"00",x"EF",x"00",x"00",x"00",x"00",x"00",x"E8",x"E8",x"E8",x"E7",x"E8",x"E8",x"E8",x"00",x"E9",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"E9",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"E9",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E8",x"E8",x"E8",x"E7",x"E8",x"E8",x"E8",x"00",x"E9",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"E9",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"E9",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"00",x"00",x"00",x"00",x"EF",x"E8",x"EF",x"EF",x"E8",x"E8",x"E8",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"EF",x"F0",x"F7",x"EF",x"00",x"EF",x"00",x"01",x"00",x"00",x"00",x"E8",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"00",x"E7",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"00",x"E7",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"00",x"E7",x"E8",x"E8",x"E8",x"E7",x"E8",x"E8",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"E8",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"00",x"E7",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"00",x"E7",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"00",x"E7",x"E8",x"E8",x"E8",x"E7",x"E8",x"E9",x"00",x"E8",x"E8",x"EF",x"EF",x"EF",x"E8",x"F7",x"EF",x"E8",x"E8",x"E8",x"01",x"EF",x"EF",x"EF",x"EF",x"00",x"00",x"01",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"EF",x"EF",x"EF",x"EF",x"00",x"EF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"E8",x"E8",x"E8",x"E8",x"F7",x"E8",x"F0",x"EF",x"E8",x"E9",x"E8",x"00",x"E9",x"E8",x"E8",x"E8",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"EF",x"EF",x"EF",x"F0",x"00",x"EF",x"00",x"00",x"01",x"00",x"00",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"E8",x"00",x"E6",x"E8",x"E7",x"E8",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E7",x"00",x"00",x"00",x"00",x"EF",x"E8",x"EF",x"F7",x"E8",x"E8",x"E8",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"EF",x"F7",x"EF",x"EF",x"00",x"00",x"00",x"00",x"00",x"00",x"E9",x"E8",x"E8",x"00",x"E9",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"E9",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"E9",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E9",x"E8",x"E8",x"00",x"E9",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"E9",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"E9",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"00",x"00",x"00",x"00",x"EE",x"E8",x"F7",x"EF",x"E7",x"E8",x"E8",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"EF",x"00",x"00",x"EF",x"00",x"00",x"00",x"00",x"00",x"00",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E9",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E9",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E9",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E9",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E9",x"E8",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E9",x"E8",x"E8",x"E8",x"00",x"E9",x"E8",x"E8",x"E8",x"00",x"00",x"00",x"00",x"EC",x"E8",x"EF",x"EF",x"E8",x"E8",x"E8",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"EF",x"00",x"EF",x"EF",x"00",x"EF",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"ED",x"E8",x"F7",x"E8",x"F5",x"E8",x"E8",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"EF",x"EF",x"EF",x"EF",x"EF",x"EF",x"00",x"00",x"00",x"00",x"00",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"E8",x"00",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"01",x"00",x"00",x"00",x"F0",x"E9",x"EF",x"E8",x"ED",x"E8",x"E8",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"EF",x"F0",x"F7",x"EF",x"00",x"EF",x"00",x"00",x"00",x"00",x"00",x"E8",x"E8",x"E8",x"E7",x"E8",x"E8",x"E8",x"00",x"E9",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"E9",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"E9",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E8",x"E8",x"E8",x"E7",x"E8",x"E8",x"E8",x"00",x"E9",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"E9",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"E9",x"E8",x"E8",x"E8",x"E8",x"E8",x"E8",x"00",x"00",x"00",x"00",x"00",x"EE",x"E8",x"F7",x"E8",x"EF",x"E8",x"E8",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"F0",x"F0",x"EF",x"EF",x"00",x"F1",x"00",x"01",x"00",x"00",x"00",x"E8",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"00",x"E7",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"00",x"E7",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"00",x"E7",x"E8",x"E8",x"E8",x"E7",x"E8",x"E8",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"E8",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"00",x"E7",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"00",x"E7",x"E8",x"E8",x"E8",x"E8",x"E7",x"E8",x"00",x"E7",x"E8",x"E8",x"E8",x"E7",x"E8",x"E9",x"00",x"E8",x"E8",x"EF",x"EF",x"F7",x"E8",x"EF",x"E8",x"F7",x"E8",x"E8",x"00",x"EF",x"EF",x"EF",x"EF",x"00",x"00",x"01",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"EF",x"ED",x"EF",x"EF",x"00",x"ED",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"E8",x"E8",x"E8",x"E8",x"EF",x"E8",x"EF",x"E8",x"EF",x"E8",x"E8",x"00",x"E9",x"E8",x"E8",x"E8",x"00",x"00",x"00",x"00")
	
	);
	
	constant bg_G : ROM :=
	(
	
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"CE",x"CE",x"CE",x"CE",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"CE",x"CE",x"CE",x"CE",x"CE",x"CE",x"CE",x"CE",x"CE",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"CE",x"CE",x"CE",x"CE",x"CE",x"CE",x"CE",x"CE",x"CE",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"CE",x"CE",x"CE",x"CE",x"CE",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"59",x"59",x"59",x"CF",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"CE",x"5A",x"59",x"59",x"5A",x"59",x"5A",x"59",x"CF",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"CE",x"5A",x"59",x"59",x"5A",x"59",x"5A",x"59",x"CF",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"CE",x"5A",x"5A",x"5A",x"5A",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"59",x"5A",x"5A",x"D6",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"CD",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"D6",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"CD",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"D6",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"CD",x"5A",x"5A",x"5A",x"5A",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"5A",x"59",x"5A",x"CE",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"CE",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"CD",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"CE",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"CD",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"CE",x"5A",x"5A",x"5A",x"5A",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"5A",x"5A",x"5A",x"D6",x"01",x"00",x"00",x"00",x"01",x"00",x"00",x"CE",x"58",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"D6",x"01",x"00",x"00",x"00",x"01",x"00",x"00",x"CE",x"58",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"D6",x"01",x"00",x"00",x"00",x"01",x"00",x"00",x"CE",x"5A",x"5A",x"5A",x"5A",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"5A",x"5A",x"5A",x"CE",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"CE",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"CE",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"CE",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"CE",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"CE",x"5A",x"5A",x"5A",x"5A",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"5A",x"5A",x"59",x"D6",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"CE",x"5A",x"59",x"5A",x"5B",x"5B",x"5B",x"59",x"D6",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"CE",x"5A",x"59",x"5A",x"5B",x"5B",x"5B",x"59",x"D6",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"CE",x"5A",x"5A",x"5A",x"5A",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"CF",x"CE",x"CE",x"CE",x"CE",x"CE",x"CE",x"CE",x"CE",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"CE",x"CE",x"CE",x"CE",x"CE",x"CE",x"CE",x"CE",x"CE",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"CE",x"CE",x"CE",x"CE",x"CE",x"CE",x"CE",x"CE",x"CE",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"5A",x"5A",x"5B",x"59",x"59",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"5A",x"5B",x"5A",x"5A",x"59",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"5A",x"5B",x"5A",x"5A",x"59",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"5A",x"59",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"5B",x"5A",x"5A",x"5A",x"5A",x"5B",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"59",x"00",x"5A",x"5A",x"5A",x"5A",x"5A",x"5B",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"59",x"00",x"5A",x"5A",x"5A",x"5A",x"5A",x"5B",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"5B",x"5A",x"5A",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"5A",x"5A",x"5A",x"01",x"5A",x"5A",x"5A",x"5A",x"59",x"5A",x"5B",x"00",x"5A",x"5A",x"5A",x"5A",x"59",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"59",x"5A",x"5B",x"00",x"5A",x"5A",x"5A",x"5A",x"59",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"59",x"5A",x"5B",x"00",x"5A",x"5A",x"5B",x"5A",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"5B",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"59",x"00",x"5A",x"5A",x"5A",x"59",x"59",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"59",x"00",x"5A",x"5A",x"5A",x"59",x"59",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"59",x"00",x"5A",x"5A",x"5A",x"5A",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"5A",x"5A",x"5A",x"5A",x"59",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"5A",x"5A",x"5A",x"5B",x"5A",x"5A",x"5A",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"5A",x"5A",x"5A",x"5B",x"5A",x"5A",x"5A",x"00",x"5B",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"5A",x"5A",x"5A",x"5B",x"5A",x"5A",x"5A",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"5A",x"5A",x"5A",x"5A",x"5B",x"5A",x"5A",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"5A",x"5A",x"5A",x"5A",x"5A",x"5B",x"5A",x"00",x"5B",x"5A",x"5A",x"5A",x"5B",x"5A",x"5A",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"5A",x"5A",x"5A",x"5A",x"5B",x"5A",x"5A",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5B",x"5A",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"59",x"5A",x"5A",x"00",x"5A",x"5A",x"5B",x"5A",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5B",x"5A",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"59",x"5A",x"5A",x"01",x"5A",x"5A",x"5A",x"5A",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"59",x"5A",x"5A",x"01",x"5B",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"59",x"5A",x"5A",x"01",x"5A",x"5A",x"5A",x"5A",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5B",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"5A",x"5A",x"5A",x"5A",x"59",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"5A",x"5A",x"5A",x"5B",x"5A",x"5A",x"5A",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"5A",x"5A",x"5A",x"5B",x"5A",x"5A",x"5A",x"00",x"5B",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"5A",x"5A",x"5A",x"5B",x"5A",x"5A",x"5A",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"5A",x"5A",x"5A",x"5A",x"5B",x"5A",x"5A",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"5A",x"5A",x"5A",x"5A",x"5A",x"5B",x"5A",x"00",x"5B",x"5A",x"5A",x"5A",x"5B",x"5A",x"5A",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"5A",x"5A",x"5A",x"5A",x"5B",x"5A",x"5A",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5B",x"5A",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"59",x"5A",x"5A",x"00",x"5A",x"5A",x"5B",x"5A",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5B",x"5A",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"59",x"5A",x"5A",x"01",x"5A",x"5A",x"5A",x"5A",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"59",x"5A",x"5A",x"01",x"5B",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"59",x"5A",x"5A",x"01",x"5A",x"5A",x"5A",x"5A",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5B",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"CE",x"CE",x"CE",x"CE",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"CE",x"CE",x"CE",x"CE",x"CE",x"CE",x"CE",x"CF",x"CE",x"5A",x"5A",x"5B",x"00",x"5A",x"5A",x"5A",x"CE",x"CE",x"CE",x"CE",x"CE",x"CE",x"CE",x"CE",x"CE",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"D6",x"CE",x"CE",x"D6",x"CE",x"CE",x"CE",x"CE",x"CE",x"5A",x"5B",x"5A",x"00",x"5A",x"5A",x"59",x"D6",x"CE",x"CE",x"D6",x"CE",x"CE",x"CE",x"CE",x"CD",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"CE",x"CE",x"CE",x"CE",x"CE",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"59",x"59",x"59",x"CF",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"CE",x"5A",x"59",x"5A",x"5A",x"59",x"5A",x"59",x"D6",x"5B",x"5A",x"5A",x"00",x"5A",x"59",x"5A",x"D6",x"5A",x"59",x"59",x"5A",x"59",x"5A",x"59",x"CF",x"5B",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"D6",x"5A",x"59",x"5A",x"5A",x"59",x"5A",x"59",x"CE",x"5B",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"CE",x"5A",x"59",x"5A",x"5A",x"59",x"5A",x"59",x"CE",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"CE",x"5A",x"5A",x"5A",x"5A",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"59",x"5A",x"5A",x"D6",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"CD",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"CE",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"D6",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"D6",x"5A",x"5B",x"5A",x"00",x"5A",x"5A",x"5A",x"CE",x"5A",x"5B",x"5A",x"5A",x"59",x"5A",x"5A",x"D6",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"D6",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"CE",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"CD",x"5A",x"5A",x"5A",x"5A",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"5A",x"59",x"5A",x"CE",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"CE",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"D6",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"CD",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"CD",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"D6",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"CE",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"CD",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"D7",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"CE",x"5A",x"5A",x"5A",x"5A",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"5A",x"5A",x"5A",x"D6",x"01",x"00",x"00",x"00",x"01",x"00",x"00",x"CE",x"59",x"5A",x"5A",x"5A",x"5B",x"5A",x"5A",x"D6",x"5A",x"5A",x"5A",x"5A",x"59",x"5A",x"5A",x"CE",x"58",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"D6",x"5A",x"5A",x"5A",x"5A",x"59",x"5A",x"5A",x"CE",x"58",x"59",x"5A",x"59",x"5A",x"5A",x"5A",x"D6",x"5A",x"5A",x"5B",x"5A",x"59",x"5A",x"5A",x"CE",x"59",x"5A",x"5A",x"5A",x"5A",x"5B",x"59",x"CE",x"01",x"00",x"00",x"00",x"01",x"00",x"00",x"CE",x"5A",x"5A",x"5A",x"5A",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"5A",x"5A",x"5A",x"CE",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"CE",x"5A",x"5A",x"5A",x"5A",x"5A",x"59",x"5A",x"CE",x"5A",x"59",x"5A",x"59",x"5A",x"5A",x"5A",x"D6",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"CE",x"5A",x"59",x"5A",x"5A",x"5B",x"5A",x"5B",x"D6",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"CE",x"5A",x"59",x"5B",x"58",x"5A",x"5A",x"5A",x"D7",x"5A",x"5A",x"59",x"5A",x"5A",x"5B",x"5A",x"D6",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"CE",x"5A",x"5A",x"5A",x"5A",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"5A",x"5A",x"59",x"D6",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"CE",x"5A",x"59",x"5A",x"5B",x"5A",x"5A",x"59",x"D6",x"5A",x"5A",x"5B",x"5A",x"5A",x"5B",x"5A",x"CE",x"5A",x"59",x"5A",x"5B",x"5B",x"5B",x"59",x"D6",x"5A",x"5A",x"5B",x"5A",x"5B",x"5A",x"5A",x"CE",x"5A",x"59",x"5A",x"5B",x"59",x"5A",x"59",x"D6",x"5A",x"5A",x"5B",x"5A",x"5A",x"5A",x"5A",x"CE",x"5A",x"59",x"5A",x"5B",x"5A",x"5A",x"59",x"CE",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"CE",x"5A",x"5A",x"5A",x"5A",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"CF",x"CE",x"CE",x"CE",x"CE",x"CE",x"CE",x"CE",x"CE",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"CE",x"D5",x"CE",x"D6",x"CE",x"D6",x"CE",x"D6",x"CE",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"CE",x"D5",x"CE",x"D6",x"CE",x"D6",x"CE",x"D6",x"CE",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"CE",x"D5",x"CE",x"D6",x"CE",x"D6",x"CE",x"D6",x"CE",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"D6",x"CE",x"CE",x"CE",x"CE",x"CE",x"CE",x"CE",x"CE",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"5A",x"5A",x"5B",x"59",x"59",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"5A",x"5B",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"5A",x"5B",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"5A",x"5B",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"5A",x"5B",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"59",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"5A",x"59",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"5A",x"59",x"5A",x"00",x"5B",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"5A",x"59",x"5A",x"00",x"5B",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"5A",x"59",x"5A",x"00",x"5B",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5B",x"5A",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"5B",x"5A",x"5A",x"5A",x"5A",x"5B",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"59",x"00",x"5A",x"5A",x"5A",x"5A",x"5A",x"5B",x"5A",x"00",x"5A",x"5A",x"5A",x"5B",x"5A",x"5A",x"59",x"00",x"5A",x"5A",x"5A",x"5A",x"5A",x"5B",x"5A",x"00",x"5A",x"5A",x"5A",x"5B",x"5A",x"5A",x"59",x"00",x"5A",x"5A",x"5A",x"5A",x"5A",x"5B",x"5A",x"00",x"5A",x"5A",x"5A",x"5B",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"59",x"5A",x"5A",x"5B",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"5B",x"5A",x"5A",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"5A",x"5A",x"5A",x"01",x"5A",x"5A",x"5A",x"5A",x"59",x"5A",x"5B",x"00",x"5A",x"5A",x"5A",x"5A",x"59",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"59",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"59",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"59",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"59",x"5A",x"5B",x"00",x"5A",x"5A",x"5B",x"5A",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"5B",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"59",x"00",x"5A",x"5A",x"5A",x"59",x"59",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"59",x"00",x"5A",x"5A",x"5A",x"59",x"59",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"59",x"00",x"5A",x"5A",x"5A",x"59",x"59",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"59",x"00",x"5A",x"5A",x"5A",x"59",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"59",x"00",x"5A",x"5A",x"5A",x"5A",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"5A",x"59",x"5A",x"5A",x"59",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"59",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"59",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"59",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"5B",x"00",x"00",x"00",x"00",x"00",x"00",x"5B",x"5A",x"5A",x"5A",x"00",x"59",x"59",x"5B",x"5A",x"59",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"59",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"59",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"5A",x"5A",x"5A",x"5B",x"5A",x"5A",x"5A",x"00",x"5B",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"5B",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"5B",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"5A",x"5B",x"5A",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"5A",x"5A",x"00",x"5A",x"5B",x"5B",x"5A",x"5A",x"5A",x"5A",x"00",x"5B",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"5B",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"5B",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"BD",x"BD",x"BD",x"BD",x"00",x"00",x"00",x"00",x"00",x"01",x"5A",x"5A",x"5A",x"5A",x"5A",x"5B",x"5A",x"00",x"5B",x"5A",x"5A",x"5A",x"5A",x"5B",x"5A",x"00",x"5B",x"5A",x"5A",x"5A",x"5A",x"5B",x"5A",x"00",x"5B",x"5A",x"5A",x"5A",x"5A",x"5B",x"5A",x"00",x"5A",x"5A",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"5A",x"00",x"59",x"5A",x"5A",x"5B",x"5A",x"5B",x"5A",x"00",x"5B",x"5A",x"5A",x"5A",x"5A",x"5B",x"5A",x"00",x"5B",x"5A",x"5A",x"5A",x"5A",x"5B",x"5A",x"00",x"5B",x"5A",x"5A",x"5A",x"5B",x"5A",x"5A",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"BD",x"BD",x"FE",x"FE",x"FE",x"FE",x"BD",x"BD",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"BD",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"BD",x"00",x"00",x"00",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"59",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"59",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"59",x"5A",x"5A",x"00",x"59",x"5B",x"5A",x"5A",x"5A",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"5A",x"5A",x"5B",x"59",x"00",x"5A",x"5A",x"5A",x"5A",x"59",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"59",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"59",x"5A",x"5A",x"00",x"5A",x"5A",x"5B",x"5A",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"BE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"BD",x"00",x"00",x"59",x"5A",x"5A",x"01",x"5B",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"5B",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"5B",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"5A",x"5A",x"5A",x"5B",x"00",x"5B",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"5B",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"5B",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"BD",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FF",x"BE",x"01",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5B",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5B",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5B",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5B",x"5B",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"5B",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5B",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5B",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5B",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"01",x"00",x"00",x"00",x"BD",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"BD",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"BE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FF",x"FE",x"BD",x"00",x"5A",x"5A",x"5A",x"5B",x"59",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"59",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"59",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"5A",x"5A",x"5A",x"5A",x"59",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"59",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"59",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"BD",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"BD",x"00",x"5A",x"5A",x"5A",x"5B",x"5A",x"5A",x"5A",x"00",x"5B",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"5B",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"5B",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"5A",x"5A",x"5A",x"5B",x"5A",x"5A",x"5A",x"00",x"5B",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"5B",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"5B",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"BD",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FD",x"FE",x"BD",x"00",x"5A",x"5A",x"5A",x"5A",x"5A",x"5B",x"5A",x"00",x"5B",x"5A",x"5A",x"5A",x"5A",x"5B",x"5A",x"00",x"5B",x"5A",x"5A",x"5A",x"5A",x"5B",x"5A",x"00",x"5B",x"5A",x"5A",x"5A",x"5B",x"5A",x"5A",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"5A",x"5A",x"5A",x"5A",x"5A",x"5B",x"5A",x"00",x"5B",x"5A",x"5A",x"5A",x"5A",x"5B",x"5A",x"00",x"5B",x"5A",x"5A",x"5A",x"5A",x"5B",x"5A",x"00",x"5B",x"5A",x"5A",x"5A",x"5B",x"5A",x"5A",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"BD",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"BD",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"01",x"00",x"00",x"BE",x"BD",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"BD",x"BC",x"00",x"00",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"59",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"59",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"59",x"5A",x"5A",x"00",x"5A",x"5A",x"5B",x"5A",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"59",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"59",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"59",x"5A",x"5A",x"00",x"5A",x"5A",x"5B",x"5A",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"BD",x"BD",x"BD",x"FE",x"FE",x"FE",x"FE",x"BD",x"BD",x"BD",x"00",x"00",x"00",x"59",x"5A",x"5A",x"01",x"5B",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"5B",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"5B",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"59",x"5A",x"5A",x"01",x"5B",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"5B",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"5B",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"BD",x"BD",x"BD",x"BD",x"BD",x"BD",x"BD",x"BD",x"00",x"00",x"01",x"01",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5B",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5B",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5B",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5B",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5B",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5B",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"BD",x"BC",x"BE",x"BD",x"BC",x"BD",x"BC",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"CE",x"D6",x"CE",x"CD",x"D6",x"CE",x"00",x"00",x"00",x"00",x"00",x"5A",x"5A",x"5A",x"5A",x"59",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"59",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"59",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"5A",x"5A",x"5A",x"5A",x"59",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"59",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"59",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"00",x"00",x"00",x"00",x"CE",x"5A",x"CF",x"CE",x"CE",x"5A",x"5A",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"CE",x"CE",x"CE",x"CD",x"00",x"CE",x"00",x"00",x"00",x"00",x"00",x"5A",x"5A",x"5A",x"5B",x"5A",x"5A",x"5A",x"00",x"5B",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"5B",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"5B",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"5A",x"5A",x"5A",x"5B",x"5A",x"5A",x"5A",x"00",x"5B",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"5B",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"5B",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"00",x"00",x"00",x"00",x"CE",x"5A",x"CE",x"CE",x"5A",x"5A",x"5A",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"CE",x"CF",x"D6",x"CE",x"00",x"CE",x"00",x"00",x"00",x"00",x"00",x"5A",x"5A",x"5A",x"5A",x"5A",x"5B",x"5A",x"00",x"5B",x"5A",x"5A",x"5A",x"5A",x"5B",x"5A",x"00",x"5B",x"5A",x"5A",x"5A",x"5A",x"5B",x"5A",x"00",x"5B",x"5A",x"5A",x"5A",x"5B",x"5A",x"5A",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"5A",x"5A",x"5A",x"5A",x"5A",x"5B",x"5A",x"00",x"5B",x"5A",x"5A",x"5A",x"5A",x"5B",x"5A",x"00",x"5B",x"5A",x"5A",x"5A",x"5A",x"5B",x"5A",x"00",x"5B",x"5A",x"5A",x"5A",x"5A",x"5A",x"59",x"00",x"5A",x"5A",x"CE",x"CE",x"CE",x"5A",x"D6",x"CE",x"5A",x"5A",x"5A",x"00",x"CE",x"CE",x"CE",x"CE",x"00",x"00",x"01",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"CE",x"CE",x"CE",x"CE",x"00",x"CE",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"5A",x"5A",x"5A",x"5A",x"D6",x"5A",x"CF",x"CE",x"5A",x"5B",x"5A",x"00",x"59",x"5A",x"5A",x"5A",x"00",x"00",x"00",x"01"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"CE",x"CE",x"CE",x"CD",x"00",x"CE",x"00",x"00",x"00",x"00",x"00",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"59",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"59",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"59",x"5A",x"5A",x"00",x"5A",x"5A",x"5B",x"5A",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"59",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"59",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"59",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5B",x"00",x"00",x"00",x"00",x"CE",x"5A",x"CE",x"D6",x"5A",x"5A",x"5A",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"CE",x"D6",x"CE",x"CE",x"00",x"00",x"00",x"00",x"00",x"00",x"59",x"5A",x"5A",x"01",x"5B",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"5B",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"5B",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"59",x"5A",x"5A",x"01",x"5B",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"5B",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"5B",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"00",x"00",x"00",x"00",x"CD",x"5A",x"D6",x"CE",x"5B",x"5A",x"5A",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"CE",x"00",x"00",x"CE",x"01",x"00",x"00",x"00",x"01",x"00",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5B",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5B",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5B",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5B",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5B",x"5A",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5B",x"5A",x"5A",x"5A",x"00",x"59",x"5A",x"5A",x"5A",x"00",x"00",x"00",x"00",x"CE",x"5A",x"CE",x"CE",x"58",x"5A",x"5A",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"CE",x"01",x"CE",x"CE",x"01",x"CE",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"CF",x"5A",x"D6",x"5A",x"D7",x"5A",x"5A",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"CE",x"CE",x"CE",x"CE",x"CE",x"CE",x"00",x"00",x"00",x"00",x"00",x"5A",x"5A",x"5A",x"5A",x"59",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"59",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"59",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"5A",x"5A",x"5A",x"5A",x"59",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"59",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"59",x"5A",x"5A",x"00",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"00",x"00",x"00",x"00",x"CF",x"5B",x"CE",x"5A",x"CF",x"5A",x"5A",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"CE",x"CD",x"D6",x"CE",x"00",x"CE",x"00",x"00",x"00",x"00",x"00",x"5A",x"5A",x"5A",x"5B",x"5A",x"5A",x"5A",x"00",x"5B",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"5B",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"5B",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"5A",x"5A",x"5A",x"5B",x"5A",x"5A",x"5A",x"00",x"5B",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"5B",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"5B",x"5A",x"5A",x"5A",x"5A",x"5A",x"5A",x"00",x"00",x"00",x"00",x"00",x"CD",x"5A",x"D6",x"5A",x"CE",x"5A",x"5A",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"CD",x"CF",x"CE",x"CE",x"00",x"CE",x"00",x"00",x"00",x"00",x"00",x"5A",x"5A",x"5A",x"5A",x"5A",x"5B",x"5A",x"00",x"5B",x"5A",x"5A",x"5A",x"5A",x"5B",x"5A",x"00",x"5B",x"5A",x"5A",x"5A",x"5A",x"5B",x"5A",x"00",x"5B",x"5A",x"5A",x"5A",x"5B",x"5A",x"5A",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"5A",x"5A",x"5A",x"5A",x"5A",x"5B",x"5A",x"00",x"5B",x"5A",x"5A",x"5A",x"5A",x"5B",x"5A",x"00",x"5B",x"5A",x"5A",x"5A",x"5A",x"5B",x"5A",x"00",x"5B",x"5A",x"5A",x"5A",x"5A",x"5A",x"59",x"00",x"5A",x"5A",x"CE",x"CE",x"D6",x"5A",x"CE",x"5A",x"D6",x"5A",x"5A",x"00",x"CE",x"CE",x"CE",x"CE",x"00",x"00",x"01",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"CE",x"CF",x"CE",x"CE",x"00",x"CE",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"5A",x"5A",x"5A",x"5A",x"CE",x"5A",x"CE",x"5A",x"CE",x"5A",x"5A",x"00",x"59",x"5A",x"5A",x"5A",x"00",x"00",x"00",x"01")
	
	);
	
	constant bg_B : ROM :=
	(
	
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"AD",x"AD",x"AD",x"AD",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"AD",x"AD",x"AD",x"AD",x"AB",x"AD",x"AD",x"AD",x"AB",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"AD",x"AD",x"AD",x"AD",x"AB",x"AD",x"AD",x"AD",x"AB",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"AD",x"AD",x"AD",x"AD",x"AD",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"02",x"00",x"00",x"10",x"10",x"10",x"AE",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"AD",x"10",x"10",x"0F",x"10",x"10",x"10",x"10",x"AE",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"AD",x"10",x"10",x"0F",x"10",x"10",x"10",x"10",x"AE",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"AD",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"B5",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"AD",x"10",x"10",x"10",x"10",x"0E",x"10",x"10",x"B5",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"AD",x"10",x"10",x"10",x"10",x"0E",x"10",x"10",x"B5",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"AD",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"0F",x"10",x"AD",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"AD",x"10",x"10",x"0E",x"10",x"10",x"10",x"10",x"AC",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"AD",x"10",x"10",x"0E",x"10",x"10",x"10",x"10",x"AC",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"AD",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"B5",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"AD",x"0F",x"10",x"10",x"10",x"10",x"10",x"10",x"B5",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"AD",x"0F",x"10",x"10",x"10",x"10",x"10",x"10",x"B5",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"AD",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"12",x"10",x"0E",x"AD",x"00",x"02",x"00",x"00",x"00",x"00",x"00",x"AD",x"10",x"10",x"10",x"12",x"10",x"10",x"10",x"AD",x"00",x"02",x"00",x"00",x"00",x"00",x"00",x"AD",x"10",x"10",x"10",x"12",x"10",x"10",x"10",x"AD",x"00",x"02",x"00",x"00",x"00",x"00",x"00",x"AD",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"B5",x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"AD",x"10",x"10",x"10",x"10",x"11",x"11",x"10",x"B3",x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"AD",x"10",x"10",x"10",x"10",x"11",x"11",x"10",x"B3",x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"AD",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"AE",x"AD",x"AD",x"AD",x"AD",x"AD",x"AD",x"AD",x"AD",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"AD",x"AD",x"AD",x"AD",x"AD",x"AD",x"AD",x"AD",x"AD",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"AD",x"AD",x"AD",x"AD",x"AD",x"AD",x"AD",x"AD",x"AD",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"0E",x"10",x"11",x"0F",x"0F",x"10",x"10",x"00",x"10",x"12",x"10",x"10",x"10",x"10",x"10",x"00",x"12",x"11",x"10",x"10",x"0F",x"10",x"10",x"00",x"10",x"12",x"10",x"10",x"10",x"10",x"10",x"00",x"12",x"11",x"10",x"10",x"0F",x"10",x"10",x"00",x"10",x"12",x"10",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"11",x"10",x"10",x"10",x"12",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"0F",x"00",x"10",x"10",x"10",x"10",x"12",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"0F",x"00",x"10",x"10",x"10",x"10",x"12",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"10",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"0F",x"10",x"11",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"0F",x"10",x"11",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"0F",x"10",x"11",x"00",x"0F",x"10",x"10",x"10",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"0E",x"10",x"10",x"10",x"0F",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"0E",x"10",x"10",x"10",x"0F",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"10",x"0F",x"10",x"10",x"00",x"10",x"12",x"10",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"02",x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"11",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"02",x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"02",x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"10",x"12",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"02",x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"00",x"0F",x"10",x"10",x"10",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"0F",x"10",x"10",x"00",x"0F",x"10",x"10",x"10",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"00",x"0F",x"10",x"10",x"10",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"02",x"12",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"02",x"12",x"10",x"10",x"00",x"11",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"02",x"12",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"00",x"10",x"10",x"10",x"11",x"10",x"10",x"10",x"02",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"10",x"0F",x"10",x"10",x"00",x"10",x"12",x"10",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"02",x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"11",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"02",x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"02",x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"10",x"12",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"02",x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"00",x"0F",x"10",x"10",x"10",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"0F",x"10",x"10",x"00",x"0F",x"10",x"10",x"10",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"00",x"0F",x"10",x"10",x"10",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"02",x"12",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"02",x"12",x"10",x"10",x"00",x"11",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"02",x"12",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"00",x"10",x"10",x"10",x"11",x"10",x"10",x"10",x"02",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"AD",x"AD",x"AD",x"AD",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"AD",x"AD",x"AD",x"AD",x"AB",x"AD",x"AD",x"AE",x"AB",x"10",x"10",x"11",x"00",x"10",x"0E",x"10",x"AD",x"AD",x"AD",x"AD",x"AB",x"AD",x"AD",x"AD",x"AB",x"10",x"10",x"10",x"00",x"10",x"0E",x"10",x"B5",x"AD",x"AD",x"B5",x"AB",x"AD",x"AD",x"AD",x"AB",x"10",x"11",x"10",x"00",x"10",x"0E",x"0F",x"B5",x"AD",x"AD",x"B5",x"AB",x"AD",x"AD",x"AD",x"AA",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"AD",x"AD",x"AD",x"AD",x"AD",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"02",x"00",x"00",x"10",x"10",x"10",x"AE",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"AD",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"B5",x"10",x"10",x"10",x"00",x"10",x"0F",x"10",x"B3",x"10",x"10",x"0F",x"10",x"10",x"10",x"10",x"AE",x"10",x"10",x"10",x"00",x"10",x"10",x"10",x"B3",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"AD",x"10",x"10",x"10",x"00",x"10",x"10",x"10",x"AB",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"AD",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"AD",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"B5",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"AD",x"10",x"10",x"10",x"10",x"0E",x"10",x"10",x"AD",x"10",x"10",x"10",x"00",x"10",x"10",x"10",x"B5",x"10",x"10",x"10",x"10",x"0E",x"10",x"10",x"B5",x"10",x"11",x"10",x"00",x"10",x"10",x"10",x"AD",x"10",x"11",x"10",x"10",x"0D",x"10",x"10",x"B5",x"10",x"10",x"10",x"00",x"10",x"10",x"10",x"B5",x"10",x"10",x"10",x"10",x"0E",x"10",x"10",x"AD",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"AD",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"0F",x"10",x"AD",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"AD",x"10",x"10",x"0E",x"10",x"10",x"10",x"10",x"B5",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"AD",x"10",x"10",x"0E",x"10",x"10",x"10",x"10",x"AC",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"B6",x"10",x"10",x"0E",x"10",x"10",x"10",x"10",x"AD",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"AD",x"10",x"10",x"0E",x"10",x"10",x"10",x"10",x"B6",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"AD",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"B5",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"AD",x"10",x"10",x"10",x"10",x"11",x"10",x"10",x"B5",x"10",x"10",x"10",x"10",x"10",x"10",x"0E",x"AD",x"0F",x"10",x"10",x"10",x"10",x"10",x"10",x"B5",x"10",x"10",x"10",x"10",x"10",x"10",x"0E",x"AD",x"0F",x"0F",x"10",x"0F",x"10",x"10",x"10",x"B5",x"10",x"10",x"11",x"10",x"10",x"10",x"0E",x"AD",x"10",x"10",x"10",x"10",x"10",x"11",x"0F",x"AD",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"AD",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"12",x"10",x"0E",x"AD",x"00",x"02",x"00",x"00",x"00",x"00",x"00",x"AD",x"10",x"10",x"10",x"12",x"10",x"0F",x"10",x"AD",x"10",x"10",x"10",x"10",x"10",x"10",x"0E",x"B5",x"10",x"10",x"10",x"12",x"10",x"10",x"10",x"AD",x"10",x"10",x"10",x"11",x"11",x"10",x"0F",x"B5",x"10",x"10",x"10",x"12",x"10",x"10",x"10",x"AD",x"10",x"10",x"11",x"0F",x"10",x"10",x"0E",x"B6",x"10",x"10",x"0F",x"12",x"10",x"11",x"10",x"B5",x"00",x"02",x"00",x"00",x"00",x"00",x"00",x"AD",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"B5",x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"AD",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"B3",x"10",x"10",x"10",x"10",x"10",x"11",x"10",x"AD",x"10",x"10",x"10",x"10",x"11",x"11",x"10",x"B3",x"10",x"10",x"10",x"10",x"11",x"10",x"10",x"AD",x"10",x"10",x"10",x"10",x"0F",x"10",x"10",x"B3",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"AD",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"AB",x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"AD",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"AE",x"AD",x"AD",x"AD",x"AD",x"AD",x"AD",x"AD",x"AD",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"AD",x"B4",x"AD",x"B5",x"AD",x"B5",x"AD",x"B5",x"AD",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"AD",x"B4",x"AD",x"B5",x"AD",x"B5",x"AD",x"B5",x"AD",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"AD",x"B4",x"AD",x"B5",x"AD",x"B5",x"AD",x"B5",x"AD",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"B5",x"AD",x"AD",x"AD",x"AD",x"AD",x"AD",x"AD",x"AD",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"0E",x"10",x"11",x"0F",x"0F",x"10",x"10",x"00",x"10",x"12",x"10",x"10",x"10",x"10",x"10",x"00",x"12",x"11",x"10",x"10",x"10",x"10",x"10",x"00",x"10",x"12",x"10",x"10",x"10",x"10",x"10",x"00",x"12",x"11",x"10",x"10",x"10",x"10",x"10",x"00",x"10",x"12",x"10",x"10",x"10",x"10",x"10",x"00",x"12",x"11",x"10",x"10",x"10",x"10",x"10",x"00",x"10",x"12",x"10",x"10",x"10",x"11",x"10",x"00",x"12",x"10",x"10",x"10",x"0F",x"10",x"10",x"00",x"10",x"12",x"10",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"10",x"0F",x"10",x"00",x"11",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"10",x"0F",x"10",x"00",x"11",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"10",x"0F",x"10",x"00",x"11",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"10",x"10",x"11",x"10",x"10",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"11",x"10",x"10",x"10",x"12",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"0F",x"00",x"10",x"10",x"10",x"10",x"12",x"10",x"10",x"00",x"10",x"10",x"10",x"11",x"10",x"10",x"0F",x"00",x"10",x"10",x"10",x"10",x"12",x"10",x"10",x"00",x"10",x"10",x"10",x"11",x"10",x"10",x"0F",x"00",x"10",x"10",x"10",x"10",x"12",x"10",x"10",x"00",x"10",x"10",x"10",x"11",x"10",x"10",x"10",x"00",x"10",x"10",x"0F",x"10",x"12",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"10",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"0F",x"10",x"11",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"0F",x"10",x"11",x"00",x"0F",x"10",x"10",x"10",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"0E",x"10",x"10",x"10",x"0F",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"0E",x"10",x"10",x"10",x"0F",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"0E",x"10",x"10",x"10",x"0F",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"0E",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"0F",x"10",x"10",x"0F",x"10",x"10",x"00",x"10",x"12",x"10",x"10",x"0F",x"10",x"10",x"00",x"10",x"12",x"10",x"10",x"0F",x"10",x"10",x"00",x"10",x"12",x"10",x"10",x"10",x"10",x"10",x"02",x"10",x"10",x"12",x"10",x"11",x"00",x"00",x"02",x"02",x"00",x"00",x"11",x"10",x"10",x"10",x"00",x"0F",x"10",x"11",x"10",x"0F",x"10",x"10",x"00",x"10",x"12",x"10",x"10",x"0F",x"10",x"10",x"00",x"10",x"12",x"10",x"10",x"0F",x"10",x"10",x"00",x"10",x"12",x"10",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"11",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"11",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"11",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"11",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"11",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"11",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"BD",x"BD",x"BD",x"BD",x"00",x"00",x"00",x"00",x"00",x"01",x"10",x"10",x"10",x"10",x"12",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"12",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"12",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"10",x"10",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"00",x"11",x"10",x"10",x"11",x"12",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"12",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"12",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"BD",x"BD",x"FE",x"FE",x"FE",x"FE",x"BD",x"BD",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"BD",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"BD",x"00",x"00",x"00",x"10",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"0F",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"0F",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"0F",x"10",x"10",x"00",x"0F",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"10",x"11",x"10",x"00",x"10",x"10",x"10",x"10",x"0F",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"0F",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"0F",x"10",x"10",x"00",x"0F",x"10",x"10",x"10",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"BE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"BD",x"00",x"02",x"12",x"10",x"10",x"00",x"11",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"11",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"11",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"02",x"00",x"00",x"10",x"10",x"10",x"11",x"00",x"11",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"11",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"11",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"BD",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FC",x"FF",x"BD",x"01",x"10",x"10",x"10",x"00",x"10",x"10",x"10",x"11",x"10",x"10",x"10",x"02",x"10",x"10",x"10",x"11",x"10",x"10",x"10",x"02",x"10",x"10",x"10",x"11",x"10",x"10",x"10",x"02",x"10",x"10",x"10",x"11",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"12",x"10",x"00",x"10",x"10",x"10",x"11",x"10",x"10",x"10",x"02",x"10",x"10",x"10",x"11",x"10",x"10",x"10",x"02",x"10",x"10",x"10",x"11",x"10",x"10",x"10",x"02",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"01",x"00",x"00",x"00",x"BD",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"BD",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"BE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FF",x"FE",x"BD",x"00",x"10",x"10",x"10",x"11",x"0F",x"10",x"10",x"00",x"10",x"12",x"10",x"10",x"0F",x"10",x"10",x"00",x"10",x"12",x"10",x"10",x"0F",x"10",x"10",x"00",x"10",x"12",x"10",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"10",x"0F",x"10",x"10",x"00",x"10",x"12",x"10",x"10",x"0F",x"10",x"10",x"00",x"10",x"12",x"10",x"10",x"0F",x"10",x"10",x"00",x"10",x"12",x"10",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"BD",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"BD",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"11",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"11",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"11",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"11",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"11",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"11",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"BD",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"BD",x"00",x"10",x"10",x"10",x"10",x"12",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"12",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"12",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"10",x"12",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"12",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"12",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"BD",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"BD",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"01",x"00",x"00",x"BE",x"BD",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"BD",x"BD",x"00",x"00",x"10",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"0F",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"0F",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"0F",x"10",x"10",x"00",x"0F",x"10",x"10",x"10",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"0F",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"0F",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"0F",x"10",x"10",x"00",x"0F",x"10",x"10",x"10",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"BD",x"BD",x"BD",x"FE",x"FE",x"FE",x"FE",x"BD",x"BD",x"BD",x"00",x"00",x"02",x"12",x"10",x"10",x"00",x"11",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"11",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"11",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"02",x"12",x"10",x"10",x"00",x"11",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"11",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"11",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"BD",x"BD",x"BD",x"BD",x"BD",x"BD",x"BD",x"BD",x"00",x"00",x"00",x"01",x"10",x"10",x"10",x"00",x"10",x"10",x"10",x"11",x"10",x"10",x"10",x"02",x"10",x"10",x"10",x"11",x"10",x"10",x"10",x"02",x"10",x"10",x"10",x"11",x"10",x"10",x"10",x"02",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"00",x"10",x"10",x"10",x"11",x"10",x"10",x"10",x"02",x"10",x"10",x"10",x"11",x"10",x"10",x"10",x"02",x"10",x"10",x"10",x"11",x"10",x"10",x"10",x"02",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"BD",x"BD",x"BD",x"BD",x"BC",x"BE",x"BD",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"AD",x"B5",x"AD",x"AD",x"B5",x"AB",x"00",x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"10",x"0F",x"10",x"10",x"00",x"10",x"12",x"10",x"10",x"0F",x"10",x"10",x"00",x"10",x"12",x"10",x"10",x"0F",x"10",x"10",x"00",x"10",x"12",x"10",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"10",x"0F",x"10",x"10",x"00",x"10",x"12",x"10",x"10",x"0F",x"10",x"10",x"00",x"10",x"12",x"10",x"10",x"0F",x"10",x"10",x"00",x"10",x"12",x"10",x"10",x"10",x"0E",x"10",x"00",x"00",x"00",x"00",x"00",x"AB",x"10",x"AD",x"AD",x"AD",x"10",x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"02",x"AD",x"AD",x"AD",x"AD",x"00",x"AD",x"00",x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"11",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"11",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"11",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"11",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"11",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"11",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"00",x"AD",x"10",x"AD",x"AD",x"10",x"12",x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"AD",x"AE",x"B5",x"AD",x"00",x"AD",x"00",x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"10",x"12",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"12",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"12",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"10",x"12",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"12",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"12",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"12",x"10",x"10",x"00",x"10",x"10",x"AD",x"AD",x"AD",x"10",x"B5",x"AD",x"10",x"10",x"10",x"00",x"AD",x"AD",x"AD",x"AD",x"00",x"00",x"01",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"AD",x"AD",x"AF",x"AD",x"00",x"AD",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"10",x"10",x"12",x"10",x"B5",x"10",x"AE",x"AD",x"10",x"11",x"10",x"00",x"10",x"10",x"10",x"0E",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"AD",x"AD",x"AD",x"AD",x"00",x"AD",x"00",x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"0F",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"0F",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"0F",x"10",x"10",x"00",x"0F",x"10",x"10",x"10",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"0F",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"0F",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"0F",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"AD",x"10",x"AD",x"B5",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"AD",x"B5",x"AD",x"AD",x"00",x"00",x"00",x"00",x"00",x"02",x"12",x"10",x"10",x"00",x"11",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"11",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"11",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"02",x"12",x"10",x"10",x"00",x"11",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"11",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"11",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"AC",x"10",x"B5",x"AD",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"AD",x"00",x"00",x"AD",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"00",x"10",x"10",x"10",x"11",x"10",x"10",x"10",x"02",x"10",x"10",x"10",x"11",x"10",x"10",x"10",x"02",x"10",x"10",x"10",x"11",x"10",x"10",x"10",x"02",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"00",x"10",x"10",x"10",x"11",x"10",x"10",x"10",x"02",x"10",x"10",x"10",x"11",x"10",x"10",x"10",x"02",x"10",x"10",x"10",x"11",x"10",x"10",x"10",x"02",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"AC",x"0E",x"AD",x"AD",x"0F",x"10",x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"AD",x"00",x"AD",x"AD",x"00",x"AD",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"02",x"00",x"00",x"00",x"AD",x"10",x"B5",x"10",x"B5",x"10",x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"AD",x"AD",x"AD",x"AD",x"AD",x"AD",x"00",x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"10",x"0F",x"10",x"10",x"00",x"10",x"12",x"10",x"10",x"0F",x"10",x"10",x"00",x"10",x"12",x"10",x"10",x"0F",x"10",x"10",x"00",x"10",x"12",x"10",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"10",x"0F",x"10",x"10",x"00",x"10",x"12",x"10",x"10",x"0F",x"10",x"10",x"00",x"10",x"12",x"10",x"10",x"0F",x"10",x"10",x"00",x"10",x"12",x"10",x"10",x"10",x"0E",x"10",x"00",x"00",x"00",x"00",x"00",x"AC",x"11",x"AD",x"10",x"AD",x"10",x"12",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"AD",x"AD",x"B5",x"AD",x"00",x"AB",x"00",x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"11",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"11",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"11",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"11",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"11",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"11",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"00",x"AE",x"10",x"B5",x"10",x"AF",x"10",x"10",x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"AD",x"AE",x"AD",x"AD",x"00",x"AE",x"00",x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"10",x"12",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"12",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"12",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"10",x"12",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"12",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"12",x"10",x"10",x"00",x"10",x"10",x"10",x"10",x"12",x"10",x"10",x"00",x"10",x"10",x"AD",x"AD",x"B5",x"10",x"AD",x"10",x"B5",x"10",x"10",x"00",x"AD",x"AD",x"AD",x"AD",x"00",x"00",x"01",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"AD",x"AD",x"AD",x"AD",x"00",x"AF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"10",x"10",x"12",x"10",x"AD",x"10",x"AD",x"10",x"AF",x"10",x"10",x"00",x"10",x"10",x"10",x"0E",x"00",x"00",x"00",x"00")
	
	);
	
begin

	dat_R <= bg_R( dir_y )( dir_x );
	dat_G <= bg_G( dir_y )( dir_x );
	dat_B <= bg_B( dir_y )( dir_x );

end comp;