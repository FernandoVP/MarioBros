library ieee;

use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity start_ROM is

	Port(
	
		dir_y : in integer;
		dir_x : in integer;
		
		dat_R : out std_logic_vector( 7 downto 0 );
		dat_G : out std_logic_vector( 7 downto 0 );
		dat_B : out std_logic_vector( 7 downto 0 )
		
	);

end start_ROM;

architecture comp of start_ROM is

	type arreglo is array( 0 to 48 ) of std_logic_vector( 0 to 7 );

	type ROM is array( 0 to 28 ) of arreglo;

	constant start_R : ROM :=
	(
	
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"01",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"36",x"6E",x"59",x"03",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"28",x"6B",x"61",x"0C",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"91",x"FF",x"F0",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"6D",x"FF",x"FF",x"1F",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"8D",x"FF",x"E8",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"68",x"FF",x"FD",x"1E",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"82",x"FF",x"E3",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"5D",x"FF",x"FA",x"0F",x"00",x"00"),
		(x"00",x"00",x"0A",x"1F",x"2D",x"32",x"32",x"2C",x"1D",x"09",x"00",x"19",x"A6",x"FF",x"EA",x"3B",x"30",x"38",x"24",x"00",x"00",x"06",x"18",x"2A",x"32",x"32",x"2B",x"15",x"03",x"00",x"00",x"00",x"00",x"14",x"39",x"34",x"04",x"0D",x"25",x"32",x"33",x"04",x"12",x"8B",x"FF",x"FB",x"4C",x"2B",x"37"),
		(x"00",x"00",x"3D",x"9B",x"D8",x"EE",x"F1",x"D6",x"93",x"39",x"00",x"C0",x"FE",x"FF",x"FE",x"FA",x"FA",x"FF",x"A9",x"00",x"01",x"2C",x"7F",x"CA",x"EF",x"F1",x"D0",x"74",x"1E",x"00",x"00",x"00",x"00",x"5D",x"FF",x"F9",x"20",x"4A",x"B7",x"F0",x"F4",x"12",x"97",x"FF",x"FF",x"FF",x"FA",x"FA",x"FF"),
		(x"00",x"4A",x"AC",x"F2",x"FF",x"FF",x"FF",x"FF",x"FA",x"BE",x"00",x"D9",x"FF",x"FC",x"FF",x"FF",x"FF",x"FF",x"C0",x"00",x"00",x"A7",x"F5",x"FF",x"FF",x"FF",x"FF",x"E7",x"86",x"0D",x"00",x"00",x"00",x"61",x"FF",x"FF",x"86",x"BD",x"FF",x"FF",x"FE",x"14",x"AE",x"FF",x"FD",x"FF",x"FF",x"FF",x"FF"),
		(x"00",x"91",x"F8",x"FF",x"C7",x"A7",x"A2",x"AE",x"D9",x"E2",x"05",x"73",x"DF",x"FF",x"F6",x"A7",x"A3",x"AF",x"6F",x"00",x"00",x"CB",x"E4",x"B1",x"A8",x"B1",x"E1",x"FF",x"D1",x"45",x"00",x"00",x"00",x"5F",x"FF",x"FF",x"D9",x"CC",x"BC",x"A9",x"A2",x"0C",x"5D",x"D4",x"FF",x"FD",x"AF",x"A0",x"AC"),
		(x"00",x"B2",x"FF",x"DC",x"62",x"12",x"00",x"0C",x"54",x"96",x"07",x"00",x"86",x"FF",x"E3",x"00",x"00",x"00",x"00",x"00",x"00",x"86",x"62",x"0D",x"01",x"13",x"82",x"E5",x"F1",x"91",x"00",x"00",x"00",x"5F",x"FF",x"FE",x"EC",x"7B",x"1B",x"00",x"00",x"00",x"00",x"61",x"FF",x"FA",x"15",x"00",x"00"),
		(x"00",x"AA",x"FF",x"EB",x"9A",x"68",x"35",x"07",x"00",x"15",x"01",x"00",x"89",x"FF",x"E5",x"04",x"00",x"00",x"00",x"00",x"00",x"10",x"03",x"00",x"00",x"00",x"03",x"A8",x"FF",x"B8",x"01",x"00",x"00",x"5F",x"FF",x"FE",x"86",x"26",x"00",x"00",x"00",x"00",x"00",x"65",x"FF",x"FA",x"1B",x"00",x"00"),
		(x"00",x"61",x"D2",x"FF",x"E7",x"D2",x"B4",x"8C",x"4B",x"00",x"00",x"00",x"8A",x"FF",x"E5",x"08",x"00",x"00",x"00",x"00",x"01",x"1C",x"4D",x"72",x"7F",x"82",x"7D",x"CF",x"FF",x"CD",x"02",x"00",x"00",x"5F",x"FE",x"FE",x"49",x"01",x"00",x"00",x"00",x"00",x"00",x"68",x"FF",x"FA",x"1E",x"00",x"00"),
		(x"00",x"16",x"76",x"D2",x"E7",x"F5",x"FF",x"FF",x"C1",x"3D",x"02",x"00",x"8B",x"FF",x"E5",x"08",x"00",x"00",x"00",x"01",x"17",x"78",x"C8",x"FA",x"FF",x"FF",x"FF",x"FF",x"FF",x"D7",x"02",x"00",x"00",x"5F",x"FF",x"FE",x"2D",x"00",x"00",x"00",x"00",x"00",x"00",x"68",x"FF",x"FA",x"1F",x"00",x"00"),
		(x"00",x"00",x"05",x"21",x"5A",x"90",x"D8",x"FE",x"F3",x"A7",x"07",x"00",x"8B",x"FF",x"E6",x"08",x"00",x"00",x"00",x"0D",x"81",x"E6",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"DB",x"01",x"00",x"00",x"5F",x"FF",x"FE",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"68",x"FF",x"FA",x"1E",x"00",x"00"),
		(x"00",x"00",x"00",x"01",x"12",x"25",x"3C",x"B2",x"FF",x"D4",x"09",x"00",x"8B",x"FF",x"E5",x"05",x"00",x"00",x"00",x"17",x"CE",x"FF",x"C8",x"7A",x"5A",x"50",x"45",x"B9",x"FF",x"DB",x"01",x"00",x"00",x"5F",x"FF",x"FE",x"24",x"00",x"00",x"00",x"00",x"00",x"01",x"68",x"FF",x"FA",x"1B",x"00",x"00"),
		(x"00",x"2E",x"28",x"04",x"00",x"00",x"02",x"97",x"FF",x"E6",x"0A",x"00",x"88",x"FF",x"E8",x"19",x"00",x"00",x"00",x"1B",x"F0",x"FF",x"99",x"1B",x"00",x"00",x"19",x"B0",x"FF",x"DB",x"02",x"00",x"00",x"5F",x"FF",x"FF",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"66",x"FF",x"FA",x"2F",x"00",x"00"),
		(x"00",x"97",x"95",x"36",x"12",x"13",x"51",x"C1",x"FF",x"DD",x"0A",x"01",x"7D",x"FF",x"EF",x"58",x"16",x"09",x"00",x"19",x"E5",x"FF",x"A3",x"31",x"0F",x"2A",x"94",x"E6",x"FF",x"DB",x"01",x"00",x"00",x"5F",x"FF",x"FE",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"5E",x"FF",x"FC",x"69",x"1B",x"07"),
		(x"00",x"C3",x"FF",x"E0",x"D6",x"D6",x"E3",x"FF",x"FB",x"A9",x"07",x"00",x"63",x"E3",x"FF",x"E3",x"D6",x"E2",x"88",x"08",x"B5",x"FD",x"F5",x"DB",x"D6",x"E0",x"BE",x"E2",x"FF",x"DB",x"01",x"00",x"00",x"5F",x"FF",x"FE",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"4A",x"DA",x"FF",x"E7",x"D7",x"DF"),
		(x"00",x"79",x"D3",x"FC",x"FF",x"FF",x"FF",x"E8",x"A3",x"46",x"03",x"00",x"2B",x"8D",x"EB",x"FF",x"FF",x"FF",x"BF",x"00",x"54",x"C2",x"FF",x"FF",x"FF",x"E8",x"6A",x"C1",x"FF",x"E8",x"01",x"00",x"01",x"65",x"FF",x"FF",x"27",x"00",x"00",x"01",x"00",x"00",x"00",x"21",x"7E",x"E3",x"FF",x"FF",x"FF"),
		(x"00",x"17",x"5A",x"A2",x"C9",x"CF",x"C0",x"8D",x"3E",x"00",x"00",x"00",x"00",x"31",x"97",x"C4",x"D4",x"E6",x"92",x"00",x"02",x"68",x"B1",x"CE",x"C1",x"81",x"05",x"79",x"F1",x"B9",x"01",x"00",x"01",x"50",x"E8",x"D7",x"1F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"22",x"8E",x"C0",x"D3",x"E3"),
		(x"00",x"02",x"06",x"0A",x"0D",x"0E",x"0B",x"09",x"05",x"00",x"00",x"00",x"00",x"04",x"0A",x"0C",x"0D",x"10",x"09",x"00",x"00",x"07",x"0B",x"0D",x"0C",x"08",x"00",x"08",x"0F",x"0C",x"00",x"00",x"00",x"05",x"0F",x"0E",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"02",x"08",x"0C",x"0D",x"0F"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00")
			
	);
	
	constant start_G : ROM :=
	(
	
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"01",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"36",x"6E",x"59",x"03",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"28",x"6B",x"61",x"0C",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"91",x"FF",x"F0",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"6D",x"FF",x"FF",x"1F",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"8D",x"FF",x"E8",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"68",x"FF",x"FD",x"1E",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"82",x"FF",x"E3",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"5D",x"FF",x"FA",x"0F",x"00",x"00"),
		(x"00",x"00",x"0A",x"1F",x"2D",x"32",x"32",x"2C",x"1D",x"09",x"00",x"19",x"A6",x"FF",x"EA",x"3B",x"30",x"38",x"24",x"00",x"00",x"06",x"18",x"2A",x"32",x"32",x"2B",x"15",x"03",x"00",x"00",x"00",x"00",x"14",x"39",x"34",x"04",x"0D",x"25",x"32",x"33",x"04",x"12",x"8B",x"FF",x"FB",x"4C",x"2B",x"37"),
		(x"00",x"00",x"3D",x"9B",x"D8",x"EE",x"F1",x"D6",x"93",x"39",x"00",x"C0",x"FE",x"FF",x"FE",x"FA",x"FA",x"FF",x"A9",x"00",x"01",x"2C",x"7F",x"CA",x"EF",x"F1",x"D0",x"74",x"1E",x"00",x"00",x"00",x"00",x"5D",x"FF",x"F9",x"20",x"4A",x"B7",x"F0",x"F4",x"12",x"97",x"FF",x"FF",x"FF",x"FA",x"FA",x"FF"),
		(x"00",x"4A",x"AC",x"F2",x"FF",x"FF",x"FF",x"FF",x"FA",x"BE",x"00",x"D9",x"FF",x"FC",x"FF",x"FF",x"FF",x"FF",x"C0",x"00",x"00",x"A7",x"F5",x"FF",x"FF",x"FF",x"FF",x"E7",x"86",x"0D",x"00",x"00",x"00",x"61",x"FF",x"FF",x"86",x"BD",x"FF",x"FF",x"FE",x"14",x"AE",x"FF",x"FD",x"FF",x"FF",x"FF",x"FF"),
		(x"00",x"91",x"F8",x"FF",x"C7",x"A7",x"A2",x"AE",x"D9",x"E2",x"05",x"73",x"DF",x"FF",x"F6",x"A7",x"A3",x"AF",x"6F",x"00",x"00",x"CB",x"E4",x"B1",x"A8",x"B1",x"E1",x"FF",x"D1",x"45",x"00",x"00",x"00",x"5F",x"FF",x"FF",x"D9",x"CC",x"BC",x"A9",x"A2",x"0C",x"5D",x"D4",x"FF",x"FD",x"AF",x"A0",x"AC"),
		(x"00",x"B2",x"FF",x"DC",x"62",x"12",x"00",x"0C",x"54",x"96",x"07",x"00",x"86",x"FF",x"E3",x"00",x"00",x"00",x"00",x"00",x"00",x"86",x"62",x"0D",x"01",x"13",x"82",x"E5",x"F1",x"91",x"00",x"00",x"00",x"5F",x"FF",x"FE",x"EC",x"7B",x"1B",x"00",x"00",x"00",x"00",x"61",x"FF",x"FA",x"15",x"00",x"00"),
		(x"00",x"AA",x"FF",x"EB",x"9A",x"68",x"35",x"07",x"00",x"15",x"01",x"00",x"89",x"FF",x"E5",x"04",x"00",x"00",x"00",x"00",x"00",x"10",x"03",x"00",x"00",x"00",x"03",x"A8",x"FF",x"B8",x"01",x"00",x"00",x"5F",x"FF",x"FE",x"86",x"26",x"00",x"00",x"00",x"00",x"00",x"65",x"FF",x"FA",x"1B",x"00",x"00"),
		(x"00",x"61",x"D2",x"FF",x"E7",x"D2",x"B4",x"8C",x"4B",x"00",x"00",x"00",x"8A",x"FF",x"E5",x"08",x"00",x"00",x"00",x"00",x"01",x"1C",x"4D",x"72",x"7F",x"82",x"7D",x"CF",x"FF",x"CD",x"02",x"00",x"00",x"5F",x"FE",x"FE",x"49",x"01",x"00",x"00",x"00",x"00",x"00",x"68",x"FF",x"FA",x"1E",x"00",x"00"),
		(x"00",x"16",x"76",x"D2",x"E7",x"F5",x"FF",x"FF",x"C1",x"3D",x"02",x"00",x"8B",x"FF",x"E5",x"08",x"00",x"00",x"00",x"01",x"17",x"78",x"C8",x"FA",x"FF",x"FF",x"FF",x"FF",x"FF",x"D7",x"02",x"00",x"00",x"5F",x"FF",x"FE",x"2D",x"00",x"00",x"00",x"00",x"00",x"00",x"68",x"FF",x"FA",x"1F",x"00",x"00"),
		(x"00",x"00",x"05",x"21",x"5A",x"90",x"D8",x"FE",x"F3",x"A7",x"07",x"00",x"8B",x"FF",x"E6",x"08",x"00",x"00",x"00",x"0D",x"81",x"E6",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"DB",x"01",x"00",x"00",x"5F",x"FF",x"FE",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"68",x"FF",x"FA",x"1E",x"00",x"00"),
		(x"00",x"00",x"00",x"01",x"12",x"25",x"3C",x"B2",x"FF",x"D4",x"09",x"00",x"8B",x"FF",x"E5",x"05",x"00",x"00",x"00",x"17",x"CE",x"FF",x"C8",x"7A",x"5A",x"50",x"45",x"B9",x"FF",x"DB",x"01",x"00",x"00",x"5F",x"FF",x"FE",x"24",x"00",x"00",x"00",x"00",x"00",x"01",x"68",x"FF",x"FA",x"1B",x"00",x"00"),
		(x"00",x"2E",x"28",x"04",x"00",x"00",x"02",x"97",x"FF",x"E6",x"0A",x"00",x"88",x"FF",x"E8",x"19",x"00",x"00",x"00",x"1B",x"F0",x"FF",x"99",x"1B",x"00",x"00",x"19",x"B0",x"FF",x"DB",x"02",x"00",x"00",x"5F",x"FF",x"FF",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"66",x"FF",x"FA",x"2F",x"00",x"00"),
		(x"00",x"97",x"95",x"36",x"12",x"13",x"51",x"C1",x"FF",x"DD",x"0A",x"01",x"7D",x"FF",x"EF",x"58",x"16",x"09",x"00",x"19",x"E5",x"FF",x"A3",x"31",x"0F",x"2A",x"94",x"E6",x"FF",x"DB",x"01",x"00",x"00",x"5F",x"FF",x"FE",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"5E",x"FF",x"FC",x"69",x"1B",x"07"),
		(x"00",x"C3",x"FF",x"E0",x"D6",x"D6",x"E3",x"FF",x"FB",x"A9",x"07",x"00",x"63",x"E3",x"FF",x"E3",x"D6",x"E2",x"88",x"08",x"B5",x"FD",x"F5",x"DB",x"D6",x"E0",x"BE",x"E2",x"FF",x"DB",x"01",x"00",x"00",x"5F",x"FF",x"FE",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"4A",x"DA",x"FF",x"E7",x"D7",x"DF"),
		(x"00",x"79",x"D3",x"FC",x"FF",x"FF",x"FF",x"E8",x"A3",x"46",x"03",x"00",x"2B",x"8D",x"EB",x"FF",x"FF",x"FF",x"BF",x"00",x"54",x"C2",x"FF",x"FF",x"FF",x"E8",x"6A",x"C1",x"FF",x"E8",x"01",x"00",x"01",x"65",x"FF",x"FF",x"27",x"00",x"00",x"01",x"00",x"00",x"00",x"21",x"7E",x"E3",x"FF",x"FF",x"FF"),
		(x"00",x"17",x"5A",x"A2",x"C9",x"CF",x"C0",x"8D",x"3E",x"00",x"00",x"00",x"00",x"31",x"97",x"C4",x"D4",x"E6",x"92",x"00",x"02",x"68",x"B1",x"CE",x"C1",x"81",x"05",x"79",x"F1",x"B9",x"01",x"00",x"01",x"50",x"E8",x"D7",x"1F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"22",x"8E",x"C0",x"D3",x"E3"),
		(x"00",x"02",x"06",x"0A",x"0D",x"0E",x"0B",x"09",x"05",x"00",x"00",x"00",x"00",x"04",x"0A",x"0C",x"0D",x"10",x"09",x"00",x"00",x"07",x"0B",x"0D",x"0C",x"08",x"00",x"08",x"0F",x"0C",x"00",x"00",x"00",x"05",x"0F",x"0E",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"02",x"08",x"0C",x"0D",x"0F"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00")
	
	);
	
	constant start_B : ROM :=
	(
	
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"01",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"36",x"6E",x"59",x"03",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"28",x"6B",x"61",x"0C",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"91",x"FF",x"F0",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"6D",x"FF",x"FF",x"1F",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"8D",x"FF",x"E8",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"68",x"FF",x"FD",x"1E",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"82",x"FF",x"E3",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"5D",x"FF",x"FA",x"0F",x"00",x"00"),
		(x"00",x"00",x"0A",x"1F",x"2D",x"32",x"32",x"2C",x"1D",x"09",x"00",x"19",x"A6",x"FF",x"EA",x"3B",x"30",x"38",x"24",x"00",x"00",x"06",x"18",x"2A",x"32",x"32",x"2B",x"15",x"03",x"00",x"00",x"00",x"00",x"14",x"39",x"34",x"04",x"0D",x"25",x"32",x"33",x"04",x"12",x"8B",x"FF",x"FB",x"4C",x"2B",x"37"),
		(x"00",x"00",x"3D",x"9B",x"D8",x"EE",x"F1",x"D6",x"93",x"39",x"00",x"C0",x"FE",x"FF",x"FE",x"FA",x"FA",x"FF",x"A9",x"00",x"01",x"2C",x"7F",x"CA",x"EF",x"F1",x"D0",x"74",x"1E",x"00",x"00",x"00",x"00",x"5D",x"FF",x"F9",x"20",x"4A",x"B7",x"F0",x"F4",x"12",x"97",x"FF",x"FF",x"FF",x"FA",x"FA",x"FF"),
		(x"00",x"4A",x"AC",x"F2",x"FF",x"FF",x"FF",x"FF",x"FA",x"BE",x"00",x"D9",x"FF",x"FC",x"FF",x"FF",x"FF",x"FF",x"C0",x"00",x"00",x"A7",x"F5",x"FF",x"FF",x"FF",x"FF",x"E7",x"86",x"0D",x"00",x"00",x"00",x"61",x"FF",x"FF",x"86",x"BD",x"FF",x"FF",x"FE",x"14",x"AE",x"FF",x"FD",x"FF",x"FF",x"FF",x"FF"),
		(x"00",x"91",x"F8",x"FF",x"C7",x"A7",x"A2",x"AE",x"D9",x"E2",x"05",x"73",x"DF",x"FF",x"F6",x"A7",x"A3",x"AF",x"6F",x"00",x"00",x"CB",x"E4",x"B1",x"A8",x"B1",x"E1",x"FF",x"D1",x"45",x"00",x"00",x"00",x"5F",x"FF",x"FF",x"D9",x"CC",x"BC",x"A9",x"A2",x"0C",x"5D",x"D4",x"FF",x"FD",x"AF",x"A0",x"AC"),
		(x"00",x"B2",x"FF",x"DC",x"62",x"12",x"00",x"0C",x"54",x"96",x"07",x"00",x"86",x"FF",x"E3",x"00",x"00",x"00",x"00",x"00",x"00",x"86",x"62",x"0D",x"01",x"13",x"82",x"E5",x"F1",x"91",x"00",x"00",x"00",x"5F",x"FF",x"FE",x"EC",x"7B",x"1B",x"00",x"00",x"00",x"00",x"61",x"FF",x"FA",x"15",x"00",x"00"),
		(x"00",x"AA",x"FF",x"EB",x"9A",x"68",x"35",x"07",x"00",x"15",x"01",x"00",x"89",x"FF",x"E5",x"04",x"00",x"00",x"00",x"00",x"00",x"10",x"03",x"00",x"00",x"00",x"03",x"A8",x"FF",x"B8",x"01",x"00",x"00",x"5F",x"FF",x"FE",x"86",x"26",x"00",x"00",x"00",x"00",x"00",x"65",x"FF",x"FA",x"1B",x"00",x"00"),
		(x"00",x"61",x"D2",x"FF",x"E7",x"D2",x"B4",x"8C",x"4B",x"00",x"00",x"00",x"8A",x"FF",x"E5",x"08",x"00",x"00",x"00",x"00",x"01",x"1C",x"4D",x"72",x"7F",x"82",x"7D",x"CF",x"FF",x"CD",x"02",x"00",x"00",x"5F",x"FE",x"FE",x"49",x"01",x"00",x"00",x"00",x"00",x"00",x"68",x"FF",x"FA",x"1E",x"00",x"00"),
		(x"00",x"16",x"76",x"D2",x"E7",x"F5",x"FF",x"FF",x"C1",x"3D",x"02",x"00",x"8B",x"FF",x"E5",x"08",x"00",x"00",x"00",x"01",x"17",x"78",x"C8",x"FA",x"FF",x"FF",x"FF",x"FF",x"FF",x"D7",x"02",x"00",x"00",x"5F",x"FF",x"FE",x"2D",x"00",x"00",x"00",x"00",x"00",x"00",x"68",x"FF",x"FA",x"1F",x"00",x"00"),
		(x"00",x"00",x"05",x"21",x"5A",x"90",x"D8",x"FE",x"F3",x"A7",x"07",x"00",x"8B",x"FF",x"E6",x"08",x"00",x"00",x"00",x"0D",x"81",x"E6",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"DB",x"01",x"00",x"00",x"5F",x"FF",x"FE",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"68",x"FF",x"FA",x"1E",x"00",x"00"),
		(x"00",x"00",x"00",x"01",x"12",x"25",x"3C",x"B2",x"FF",x"D4",x"09",x"00",x"8B",x"FF",x"E5",x"05",x"00",x"00",x"00",x"17",x"CE",x"FF",x"C8",x"7A",x"5A",x"50",x"45",x"B9",x"FF",x"DB",x"01",x"00",x"00",x"5F",x"FF",x"FE",x"24",x"00",x"00",x"00",x"00",x"00",x"01",x"68",x"FF",x"FA",x"1B",x"00",x"00"),
		(x"00",x"2E",x"28",x"04",x"00",x"00",x"02",x"97",x"FF",x"E6",x"0A",x"00",x"88",x"FF",x"E8",x"19",x"00",x"00",x"00",x"1B",x"F0",x"FF",x"99",x"1B",x"00",x"00",x"19",x"B0",x"FF",x"DB",x"02",x"00",x"00",x"5F",x"FF",x"FF",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"66",x"FF",x"FA",x"2F",x"00",x"00"),
		(x"00",x"97",x"95",x"36",x"12",x"13",x"51",x"C1",x"FF",x"DD",x"0A",x"01",x"7D",x"FF",x"EF",x"58",x"16",x"09",x"00",x"19",x"E5",x"FF",x"A3",x"31",x"0F",x"2A",x"94",x"E6",x"FF",x"DB",x"01",x"00",x"00",x"5F",x"FF",x"FE",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"5E",x"FF",x"FC",x"69",x"1B",x"07"),
		(x"00",x"C3",x"FF",x"E0",x"D6",x"D6",x"E3",x"FF",x"FB",x"A9",x"07",x"00",x"63",x"E3",x"FF",x"E3",x"D6",x"E2",x"88",x"08",x"B5",x"FD",x"F5",x"DB",x"D6",x"E0",x"BE",x"E2",x"FF",x"DB",x"01",x"00",x"00",x"5F",x"FF",x"FE",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"4A",x"DA",x"FF",x"E7",x"D7",x"DF"),
		(x"00",x"79",x"D3",x"FC",x"FF",x"FF",x"FF",x"E8",x"A3",x"46",x"03",x"00",x"2B",x"8D",x"EB",x"FF",x"FF",x"FF",x"BF",x"00",x"54",x"C2",x"FF",x"FF",x"FF",x"E8",x"6A",x"C1",x"FF",x"E8",x"01",x"00",x"01",x"65",x"FF",x"FF",x"27",x"00",x"00",x"01",x"00",x"00",x"00",x"21",x"7E",x"E3",x"FF",x"FF",x"FF"),
		(x"00",x"17",x"5A",x"A2",x"C9",x"CF",x"C0",x"8D",x"3E",x"00",x"00",x"00",x"00",x"31",x"97",x"C4",x"D4",x"E6",x"92",x"00",x"02",x"68",x"B1",x"CE",x"C1",x"81",x"05",x"79",x"F1",x"B9",x"01",x"00",x"01",x"50",x"E8",x"D7",x"1F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"22",x"8E",x"C0",x"D3",x"E3"),
		(x"00",x"02",x"06",x"0A",x"0D",x"0E",x"0B",x"09",x"05",x"00",x"00",x"00",x"00",x"04",x"0A",x"0C",x"0D",x"10",x"09",x"00",x"00",x"07",x"0B",x"0D",x"0C",x"08",x"00",x"08",x"0F",x"0C",x"00",x"00",x"00",x"05",x"0F",x"0E",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"02",x"08",x"0C",x"0D",x"0F"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00")
	
	);
	
begin

	dat_R <= start_R( dir_y )( dir_x );
	dat_G <= start_G( dir_y )( dir_x );
	dat_B <= start_B( dir_y )( dir_x );

end comp;