library ieee;

use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity nivel_ROM is

	Port(
	
		dir_y : in integer;
		dir_x : in integer;
		
		dat_R : out std_logic_vector( 7 downto 0 );
		dat_G : out std_logic_vector( 7 downto 0 );
		dat_B : out std_logic_vector( 7 downto 0 )
		
	);

end nivel_ROM;

architecture comp of nivel_ROM is

	type arreglo is array( 0 to 48 ) of std_logic_vector( 0 to 7 );

	type ROM is array( 0 to 18 ) of arreglo;

	constant nivel_R : ROM :=
	(
	
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"01",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"AA",x"D2",x"36",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"62",x"D8",x"84",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"FB",x"FF",x"50",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"88",x"FF",x"B5",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"63",x"7A",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"82",x"FF",x"AE",x"00",x"00"),
		(x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"82",x"FF",x"AE",x"00",x"00"),
		(x"00",x"00",x"00",x"4D",x"65",x"17",x"15",x"47",x"59",x"4A",x"1F",x"00",x"00",x"00",x"00",x"51",x"64",x"19",x"00",x"34",x"66",x"3E",x"00",x"00",x"00",x"00",x"00",x"00",x"47",x"60",x"1F",x"00",x"00",x"01",x"26",x"48",x"56",x"58",x"4D",x"2F",x"01",x"00",x"00",x"00",x"82",x"FF",x"AE",x"00",x"00"),
		(x"00",x"00",x"00",x"E8",x"FF",x"71",x"79",x"F3",x"FF",x"F2",x"8F",x"0E",x"00",x"00",x"00",x"F2",x"FF",x"4C",x"00",x"87",x"FF",x"CA",x"12",x"00",x"00",x"00",x"00",x"11",x"E3",x"FF",x"4E",x"01",x"0A",x"4D",x"AB",x"F1",x"FF",x"FE",x"FC",x"BC",x"52",x"0A",x"00",x"01",x"81",x"FF",x"AE",x"00",x"00"),
		(x"00",x"00",x"00",x"D8",x"FF",x"D1",x"CF",x"DD",x"DF",x"FE",x"F2",x"6C",x"00",x"00",x"01",x"E1",x"FF",x"48",x"00",x"43",x"D0",x"E6",x"5D",x"00",x"00",x"00",x"00",x"69",x"F7",x"A2",x"1F",x"00",x"5F",x"E7",x"FF",x"E2",x"D5",x"D5",x"E0",x"FF",x"F7",x"4B",x"03",x"00",x"82",x"FF",x"AF",x"00",x"00"),
		(x"00",x"00",x"00",x"D9",x"FF",x"E2",x"60",x"00",x"2B",x"B4",x"FF",x"B8",x"00",x"00",x"00",x"E1",x"FF",x"48",x"00",x"0E",x"8E",x"FF",x"A2",x"00",x"00",x"00",x"00",x"C2",x"FF",x"57",x"00",x"34",x"C0",x"FF",x"A6",x"2C",x"00",x"00",x"24",x"AA",x"FF",x"B7",x"27",x"00",x"82",x"FF",x"AE",x"00",x"00"),
		(x"00",x"00",x"00",x"D8",x"FF",x"78",x"09",x"00",x"00",x"57",x"FF",x"D9",x"00",x"00",x"00",x"E1",x"FF",x"49",x"00",x"00",x"56",x"FB",x"D3",x"18",x"00",x"00",x"2F",x"F3",x"DA",x"2C",x"00",x"70",x"FC",x"BE",x"20",x"03",x"08",x"08",x"07",x"1A",x"E6",x"F8",x"3F",x"00",x"82",x"FF",x"AF",x"00",x"00"),
		(x"00",x"01",x"00",x"D8",x"FF",x"58",x"00",x"00",x"00",x"46",x"FF",x"E2",x"00",x"00",x"00",x"E1",x"FF",x"47",x"00",x"00",x"2A",x"B0",x"EF",x"66",x"00",x"02",x"90",x"FE",x"85",x"14",x"00",x"89",x"FF",x"FE",x"FC",x"FD",x"FC",x"FC",x"FC",x"FC",x"FF",x"FF",x"48",x"00",x"82",x"FF",x"AE",x"01",x"00"),
		(x"00",x"00",x"00",x"D8",x"FF",x"53",x"00",x"00",x"00",x"47",x"FF",x"E2",x"00",x"00",x"00",x"E1",x"FF",x"48",x"00",x"00",x"00",x"67",x"FE",x"B4",x"00",x"0C",x"E6",x"FF",x"36",x"00",x"00",x"8B",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FE",x"FF",x"FF",x"4D",x"00",x"82",x"FF",x"AE",x"00",x"00"),
		(x"00",x"00",x"00",x"D8",x"FF",x"53",x"01",x"00",x"00",x"47",x"FF",x"E2",x"00",x"00",x"00",x"E1",x"FF",x"48",x"00",x"00",x"00",x"3A",x"DD",x"E1",x"26",x"58",x"FC",x"C0",x"1B",x"00",x"00",x"77",x"FF",x"C0",x"2D",x"1C",x"22",x"23",x"24",x"22",x"1E",x"1A",x"07",x"00",x"82",x"FF",x"AE",x"00",x"00"),
		(x"00",x"00",x"00",x"D8",x"FF",x"53",x"00",x"00",x"00",x"47",x"FF",x"E2",x"00",x"00",x"00",x"E1",x"FF",x"48",x"00",x"00",x"00",x"16",x"8C",x"F8",x"7B",x"B8",x"FF",x"65",x"09",x"00",x"00",x"3E",x"CB",x"F9",x"91",x"28",x"00",x"00",x"00",x"03",x"30",x"8A",x"2C",x"00",x"82",x"FF",x"AE",x"00",x"00"),
		(x"00",x"01",x"00",x"D8",x"FF",x"53",x"00",x"00",x"01",x"47",x"FF",x"E2",x"00",x"00",x"00",x"E0",x"FF",x"48",x"00",x"00",x"00",x"00",x"46",x"F8",x"DD",x"F4",x"EF",x"21",x"00",x"00",x"00",x"04",x"64",x"E9",x"FF",x"D0",x"B8",x"B1",x"B1",x"BC",x"D5",x"FF",x"4D",x"00",x"82",x"FF",x"AE",x"00",x"00"),
		(x"00",x"00",x"00",x"E7",x"FF",x"59",x"00",x"00",x"00",x"4C",x"FF",x"F2",x"00",x"00",x"00",x"F1",x"FF",x"4D",x"00",x"00",x"00",x"00",x"20",x"C1",x"FF",x"FF",x"A9",x"09",x"00",x"00",x"00",x"00",x"11",x"5B",x"B1",x"EF",x"FF",x"FF",x"FF",x"FF",x"D8",x"A3",x"26",x"00",x"8B",x"FF",x"BA",x"00",x"00"),
		(x"00",x"00",x"00",x"70",x"92",x"2B",x"00",x"00",x"00",x"25",x"91",x"76",x"00",x"00",x"00",x"75",x"92",x"25",x"01",x"00",x"00",x"00",x"0A",x"46",x"88",x"84",x"39",x"04",x"00",x"00",x"00",x"01",x"00",x"00",x"28",x"5E",x"78",x"82",x"7F",x"6E",x"4A",x"16",x"01",x"00",x"44",x"95",x"5B",x"00",x"00"),
		(x"00",x"00",x"02",x"00",x"01",x"00",x"02",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"01",x"00",x"00",x"00",x"01",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00")
	
	);
	
	constant nivel_G : ROM :=
	(
	
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"01",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"AA",x"D2",x"36",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"62",x"D8",x"84",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"FB",x"FF",x"50",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"88",x"FF",x"B5",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"63",x"7A",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"82",x"FF",x"AE",x"00",x"00"),
		(x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"82",x"FF",x"AE",x"00",x"00"),
		(x"00",x"00",x"00",x"4D",x"65",x"17",x"15",x"47",x"59",x"4A",x"1F",x"00",x"00",x"00",x"00",x"51",x"64",x"19",x"00",x"34",x"66",x"3E",x"00",x"00",x"00",x"00",x"00",x"00",x"47",x"60",x"1F",x"00",x"00",x"01",x"26",x"48",x"56",x"58",x"4D",x"2F",x"01",x"00",x"00",x"00",x"82",x"FF",x"AE",x"00",x"00"),
		(x"00",x"00",x"00",x"E8",x"FF",x"71",x"79",x"F3",x"FF",x"F2",x"8F",x"0E",x"00",x"00",x"00",x"F2",x"FF",x"4C",x"00",x"87",x"FF",x"CA",x"12",x"00",x"00",x"00",x"00",x"11",x"E3",x"FF",x"4E",x"01",x"0A",x"4D",x"AB",x"F1",x"FF",x"FE",x"FC",x"BC",x"52",x"0A",x"00",x"01",x"81",x"FF",x"AE",x"00",x"00"),
		(x"00",x"00",x"00",x"D8",x"FF",x"D1",x"CF",x"DD",x"DF",x"FE",x"F2",x"6C",x"00",x"00",x"01",x"E1",x"FF",x"48",x"00",x"43",x"D0",x"E6",x"5D",x"00",x"00",x"00",x"00",x"69",x"F7",x"A2",x"1F",x"00",x"5F",x"E7",x"FF",x"E2",x"D5",x"D5",x"E0",x"FF",x"F7",x"4B",x"03",x"00",x"82",x"FF",x"AF",x"00",x"00"),
		(x"00",x"00",x"00",x"D9",x"FF",x"E2",x"60",x"00",x"2B",x"B4",x"FF",x"B8",x"00",x"00",x"00",x"E1",x"FF",x"48",x"00",x"0E",x"8E",x"FF",x"A2",x"00",x"00",x"00",x"00",x"C2",x"FF",x"57",x"00",x"34",x"C0",x"FF",x"A6",x"2C",x"00",x"00",x"24",x"AA",x"FF",x"B7",x"27",x"00",x"82",x"FF",x"AE",x"00",x"00"),
		(x"00",x"00",x"00",x"D8",x"FF",x"78",x"09",x"00",x"00",x"57",x"FF",x"D9",x"00",x"00",x"00",x"E1",x"FF",x"49",x"00",x"00",x"56",x"FB",x"D3",x"18",x"00",x"00",x"2F",x"F3",x"DA",x"2C",x"00",x"70",x"FC",x"BE",x"20",x"03",x"08",x"08",x"07",x"1A",x"E6",x"F8",x"3F",x"00",x"82",x"FF",x"AF",x"00",x"00"),
		(x"00",x"01",x"00",x"D8",x"FF",x"58",x"00",x"00",x"00",x"46",x"FF",x"E2",x"00",x"00",x"00",x"E1",x"FF",x"47",x"00",x"00",x"2A",x"B0",x"EF",x"66",x"00",x"02",x"90",x"FE",x"85",x"14",x"00",x"89",x"FF",x"FE",x"FC",x"FD",x"FC",x"FC",x"FC",x"FC",x"FF",x"FF",x"48",x"00",x"82",x"FF",x"AE",x"01",x"00"),
		(x"00",x"00",x"00",x"D8",x"FF",x"53",x"00",x"00",x"00",x"47",x"FF",x"E2",x"00",x"00",x"00",x"E1",x"FF",x"48",x"00",x"00",x"00",x"67",x"FE",x"B4",x"00",x"0C",x"E6",x"FF",x"36",x"00",x"00",x"8B",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FE",x"FF",x"FF",x"4D",x"00",x"82",x"FF",x"AE",x"00",x"00"),
		(x"00",x"00",x"00",x"D8",x"FF",x"53",x"01",x"00",x"00",x"47",x"FF",x"E2",x"00",x"00",x"00",x"E1",x"FF",x"48",x"00",x"00",x"00",x"3A",x"DD",x"E1",x"26",x"58",x"FC",x"C0",x"1B",x"00",x"00",x"77",x"FF",x"C0",x"2D",x"1C",x"22",x"23",x"24",x"22",x"1E",x"1A",x"07",x"00",x"82",x"FF",x"AE",x"00",x"00"),
		(x"00",x"00",x"00",x"D8",x"FF",x"53",x"00",x"00",x"00",x"47",x"FF",x"E2",x"00",x"00",x"00",x"E1",x"FF",x"48",x"00",x"00",x"00",x"16",x"8C",x"F8",x"7B",x"B8",x"FF",x"65",x"09",x"00",x"00",x"3E",x"CB",x"F9",x"91",x"28",x"00",x"00",x"00",x"03",x"30",x"8A",x"2C",x"00",x"82",x"FF",x"AE",x"00",x"00"),
		(x"00",x"01",x"00",x"D8",x"FF",x"53",x"00",x"00",x"01",x"47",x"FF",x"E2",x"00",x"00",x"00",x"E0",x"FF",x"48",x"00",x"00",x"00",x"00",x"46",x"F8",x"DD",x"F4",x"EF",x"21",x"00",x"00",x"00",x"04",x"64",x"E9",x"FF",x"D0",x"B8",x"B1",x"B1",x"BC",x"D5",x"FF",x"4D",x"00",x"82",x"FF",x"AE",x"00",x"00"),
		(x"00",x"00",x"00",x"E7",x"FF",x"59",x"00",x"00",x"00",x"4C",x"FF",x"F2",x"00",x"00",x"00",x"F1",x"FF",x"4D",x"00",x"00",x"00",x"00",x"20",x"C1",x"FF",x"FF",x"A9",x"09",x"00",x"00",x"00",x"00",x"11",x"5B",x"B1",x"EF",x"FF",x"FF",x"FF",x"FF",x"D8",x"A3",x"26",x"00",x"8B",x"FF",x"BA",x"00",x"00"),
		(x"00",x"00",x"00",x"70",x"92",x"2B",x"00",x"00",x"00",x"25",x"91",x"76",x"00",x"00",x"00",x"75",x"92",x"25",x"01",x"00",x"00",x"00",x"0A",x"46",x"88",x"84",x"39",x"04",x"00",x"00",x"00",x"01",x"00",x"00",x"28",x"5E",x"78",x"82",x"7F",x"6E",x"4A",x"16",x"01",x"00",x"44",x"95",x"5B",x"00",x"00"),
		(x"00",x"00",x"02",x"00",x"01",x"00",x"02",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"01",x"00",x"00",x"00",x"01",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00")
	
	);
	
	constant nivel_B : ROM :=
	(
	
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"01",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"AA",x"D2",x"36",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"62",x"D8",x"84",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"FB",x"FF",x"50",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"88",x"FF",x"B5",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"63",x"7A",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"82",x"FF",x"AE",x"00",x"00"),
		(x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"82",x"FF",x"AE",x"00",x"00"),
		(x"00",x"00",x"00",x"4D",x"65",x"17",x"15",x"47",x"59",x"4A",x"1F",x"00",x"00",x"00",x"00",x"51",x"64",x"19",x"00",x"34",x"66",x"3E",x"00",x"00",x"00",x"00",x"00",x"00",x"47",x"60",x"1F",x"00",x"00",x"01",x"26",x"48",x"56",x"58",x"4D",x"2F",x"01",x"00",x"00",x"00",x"82",x"FF",x"AE",x"00",x"00"),
		(x"00",x"00",x"00",x"E8",x"FF",x"71",x"79",x"F3",x"FF",x"F2",x"8F",x"0E",x"00",x"00",x"00",x"F2",x"FF",x"4C",x"00",x"87",x"FF",x"CA",x"12",x"00",x"00",x"00",x"00",x"11",x"E3",x"FF",x"4E",x"01",x"0A",x"4D",x"AB",x"F1",x"FF",x"FE",x"FC",x"BC",x"52",x"0A",x"00",x"01",x"81",x"FF",x"AE",x"00",x"00"),
		(x"00",x"00",x"00",x"D8",x"FF",x"D1",x"CF",x"DD",x"DF",x"FE",x"F2",x"6C",x"00",x"00",x"01",x"E1",x"FF",x"48",x"00",x"43",x"D0",x"E6",x"5D",x"00",x"00",x"00",x"00",x"69",x"F7",x"A2",x"1F",x"00",x"5F",x"E7",x"FF",x"E2",x"D5",x"D5",x"E0",x"FF",x"F7",x"4B",x"03",x"00",x"82",x"FF",x"AF",x"00",x"00"),
		(x"00",x"00",x"00",x"D9",x"FF",x"E2",x"60",x"00",x"2B",x"B4",x"FF",x"B8",x"00",x"00",x"00",x"E1",x"FF",x"48",x"00",x"0E",x"8E",x"FF",x"A2",x"00",x"00",x"00",x"00",x"C2",x"FF",x"57",x"00",x"34",x"C0",x"FF",x"A6",x"2C",x"00",x"00",x"24",x"AA",x"FF",x"B7",x"27",x"00",x"82",x"FF",x"AE",x"00",x"00"),
		(x"00",x"00",x"00",x"D8",x"FF",x"78",x"09",x"00",x"00",x"57",x"FF",x"D9",x"00",x"00",x"00",x"E1",x"FF",x"49",x"00",x"00",x"56",x"FB",x"D3",x"18",x"00",x"00",x"2F",x"F3",x"DA",x"2C",x"00",x"70",x"FC",x"BE",x"20",x"03",x"08",x"08",x"07",x"1A",x"E6",x"F8",x"3F",x"00",x"82",x"FF",x"AF",x"00",x"00"),
		(x"00",x"01",x"00",x"D8",x"FF",x"58",x"00",x"00",x"00",x"46",x"FF",x"E2",x"00",x"00",x"00",x"E1",x"FF",x"47",x"00",x"00",x"2A",x"B0",x"EF",x"66",x"00",x"02",x"90",x"FE",x"85",x"14",x"00",x"89",x"FF",x"FE",x"FC",x"FD",x"FC",x"FC",x"FC",x"FC",x"FF",x"FF",x"48",x"00",x"82",x"FF",x"AE",x"01",x"00"),
		(x"00",x"00",x"00",x"D8",x"FF",x"53",x"00",x"00",x"00",x"47",x"FF",x"E2",x"00",x"00",x"00",x"E1",x"FF",x"48",x"00",x"00",x"00",x"67",x"FE",x"B4",x"00",x"0C",x"E6",x"FF",x"36",x"00",x"00",x"8B",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FE",x"FF",x"FF",x"4D",x"00",x"82",x"FF",x"AE",x"00",x"00"),
		(x"00",x"00",x"00",x"D8",x"FF",x"53",x"01",x"00",x"00",x"47",x"FF",x"E2",x"00",x"00",x"00",x"E1",x"FF",x"48",x"00",x"00",x"00",x"3A",x"DD",x"E1",x"26",x"58",x"FC",x"C0",x"1B",x"00",x"00",x"77",x"FF",x"C0",x"2D",x"1C",x"22",x"23",x"24",x"22",x"1E",x"1A",x"07",x"00",x"82",x"FF",x"AE",x"00",x"00"),
		(x"00",x"00",x"00",x"D8",x"FF",x"53",x"00",x"00",x"00",x"47",x"FF",x"E2",x"00",x"00",x"00",x"E1",x"FF",x"48",x"00",x"00",x"00",x"16",x"8C",x"F8",x"7B",x"B8",x"FF",x"65",x"09",x"00",x"00",x"3E",x"CB",x"F9",x"91",x"28",x"00",x"00",x"00",x"03",x"30",x"8A",x"2C",x"00",x"82",x"FF",x"AE",x"00",x"00"),
		(x"00",x"01",x"00",x"D8",x"FF",x"53",x"00",x"00",x"01",x"47",x"FF",x"E2",x"00",x"00",x"00",x"E0",x"FF",x"48",x"00",x"00",x"00",x"00",x"46",x"F8",x"DD",x"F4",x"EF",x"21",x"00",x"00",x"00",x"04",x"64",x"E9",x"FF",x"D0",x"B8",x"B1",x"B1",x"BC",x"D5",x"FF",x"4D",x"00",x"82",x"FF",x"AE",x"00",x"00"),
		(x"00",x"00",x"00",x"E7",x"FF",x"59",x"00",x"00",x"00",x"4C",x"FF",x"F2",x"00",x"00",x"00",x"F1",x"FF",x"4D",x"00",x"00",x"00",x"00",x"20",x"C1",x"FF",x"FF",x"A9",x"09",x"00",x"00",x"00",x"00",x"11",x"5B",x"B1",x"EF",x"FF",x"FF",x"FF",x"FF",x"D8",x"A3",x"26",x"00",x"8B",x"FF",x"BA",x"00",x"00"),
		(x"00",x"00",x"00",x"70",x"92",x"2B",x"00",x"00",x"00",x"25",x"91",x"76",x"00",x"00",x"00",x"75",x"92",x"25",x"01",x"00",x"00",x"00",x"0A",x"46",x"88",x"84",x"39",x"04",x"00",x"00",x"00",x"01",x"00",x"00",x"28",x"5E",x"78",x"82",x"7F",x"6E",x"4A",x"16",x"01",x"00",x"44",x"95",x"5B",x"00",x"00"),
		(x"00",x"00",x"02",x"00",x"01",x"00",x"02",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"01",x"00",x"00",x"00",x"01",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00")
	
	);
	
begin

	dat_R <= nivel_R( dir_y )( dir_x );
	dat_G <= nivel_G( dir_y )( dir_x );
	dat_B <= nivel_B( dir_y )( dir_x );

end comp;