library ieee;

use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity fuego_ROM is

	Port(
	
		dir_y : in integer;
		dir_x : in integer;
		
		dat_R : out std_logic_vector( 7 downto 0 );
		dat_G : out std_logic_vector( 7 downto 0 );
		dat_B : out std_logic_vector( 7 downto 0 )
		
	);

end fuego_ROM;

architecture comp of fuego_ROM is

	type arreglo is array( 0 to 24 ) of std_logic_vector( 0 to 7 );

	type ROM is array( 0 to 8 ) of arreglo;

	constant fuego_R : ROM :=
	(
	
		(x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"F9",x"00",x"00",x"F9",x"F9",x"00",x"F9",x"FA",x"F9",x"00",x"01",x"F9",x"F9",x"00",x"00",x"00",x"00",x"01"),
		(x"00",x"00",x"00",x"00",x"01",x"F9",x"F7",x"F9",x"F9",x"F9",x"F9",x"00",x"F9",x"F9",x"F9",x"F9",x"F9",x"F8",x"F9",x"F9",x"F9",x"00",x"01",x"00",x"00"),
		(x"00",x"00",x"F9",x"F9",x"F9",x"FA",x"FF",x"FF",x"FF",x"F9",x"F7",x"F9",x"F7",x"F9",x"F9",x"F9",x"F9",x"F9",x"F9",x"F9",x"F9",x"F9",x"00",x"00",x"00"),
		(x"00",x"F9",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F9",x"F9",x"F9",x"F9",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"F9",x"F9",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FE",x"FF",x"FF",x"FA",x"F9",x"F9",x"FA",x"F9",x"F9",x"F7",x"F9",x"F9",x"FA",x"F9",x"F9",x"FC"),
		(x"00",x"F9",x"F9",x"FF",x"FE",x"FF",x"FF",x"F9",x"F9",x"FF",x"FF",x"FF",x"FF",x"FB",x"F9",x"FF",x"FF",x"F9",x"FA",x"FA",x"F9",x"F9",x"01",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"F9",x"F9",x"F9",x"FA",x"F9",x"F9",x"F9",x"F8",x"F9",x"F9",x"F9",x"F9",x"F9",x"F8",x"F9",x"F9",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"01",x"FC",x"00",x"00",x"F9",x"F9",x"F9",x"F9",x"F9",x"F9",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00")
	
	);
	
	constant fuego_G : ROM :=
	(
	
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"38",x"00",x"00",x"38",x"38",x"00",x"38",x"37",x"38",x"00",x"01",x"38",x"38",x"00",x"00",x"01",x"00",x"00"),
		(x"00",x"00",x"01",x"00",x"00",x"38",x"38",x"38",x"38",x"38",x"38",x"00",x"38",x"38",x"38",x"38",x"38",x"37",x"38",x"38",x"38",x"00",x"01",x"00",x"00"),
		(x"00",x"00",x"38",x"38",x"38",x"37",x"A0",x"A0",x"A0",x"38",x"38",x"38",x"38",x"38",x"38",x"38",x"38",x"38",x"38",x"38",x"38",x"38",x"00",x"00",x"00"),
		(x"00",x"38",x"FF",x"A0",x"A0",x"A0",x"A0",x"A1",x"A0",x"9F",x"A0",x"A0",x"A0",x"A0",x"A1",x"A0",x"38",x"38",x"38",x"38",x"00",x"01",x"00",x"00",x"00"),
		(x"00",x"38",x"38",x"FF",x"FF",x"FF",x"FF",x"A0",x"A0",x"9F",x"A0",x"A0",x"37",x"38",x"38",x"37",x"38",x"38",x"38",x"38",x"38",x"37",x"38",x"38",x"37"),
		(x"00",x"38",x"38",x"A0",x"A1",x"A1",x"A0",x"38",x"38",x"A0",x"A0",x"A0",x"A0",x"37",x"38",x"A0",x"A0",x"38",x"39",x"39",x"38",x"38",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"38",x"38",x"38",x"39",x"38",x"38",x"38",x"37",x"38",x"38",x"38",x"38",x"38",x"37",x"38",x"38",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"37",x"00",x"00",x"38",x"38",x"38",x"38",x"38",x"38",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00")
		
	);
	
	constant fuego_B : ROM :=
	(
	
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"02",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"01",x"01",x"00",x"01",x"01",x"00",x"00",x"01",x"01",x"00",x"02",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"01",x"01",x"01",x"01",x"01",x"00",x"00",x"01",x"01",x"01",x"01",x"01",x"00",x"01",x"01",x"01",x"00",x"01",x"00",x"00"),
		(x"00",x"00",x"01",x"01",x"01",x"01",x"44",x"44",x"44",x"01",x"01",x"01",x"01",x"01",x"00",x"01",x"01",x"01",x"01",x"01",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"01",x"FD",x"44",x"44",x"44",x"42",x"45",x"44",x"44",x"44",x"44",x"44",x"44",x"45",x"44",x"01",x"01",x"01",x"01",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"01",x"01",x"FF",x"FF",x"FF",x"FF",x"44",x"44",x"43",x"44",x"44",x"01",x"01",x"00",x"01",x"00",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00"),
		(x"00",x"01",x"01",x"44",x"44",x"45",x"42",x"01",x"01",x"44",x"44",x"44",x"44",x"03",x"01",x"44",x"44",x"01",x"00",x"02",x"01",x"01",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"01",x"01",x"01",x"02",x"01",x"01",x"01",x"00",x"01",x"01",x"01",x"00",x"01",x"00",x"01",x"01",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00")
		
	);
	
begin

	dat_R <= fuego_R( dir_y )( dir_x );
	dat_G <= fuego_G( dir_y )( dir_x );
	dat_B <= fuego_B( dir_y )( dir_x );

end comp;