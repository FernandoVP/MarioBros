library ieee;

use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity bloque_ROM is

	Port(
	
		dir_y : in integer;
		dir_x : in integer;
		
		dat_R : out std_logic_vector( 7 downto 0 );
		dat_G : out std_logic_vector( 7 downto 0 );
		dat_B : out std_logic_vector( 7 downto 0 )
		
	);

end bloque_ROM;

architecture comp of bloque_ROM is

	type arreglo is array( 0 to 14 ) of std_logic_vector( 0 to 7 );

	type ROM is array( 0 to 13 ) of arreglo;

	constant bloque_R : ROM :=
	(
	
		(x"FF",x"D5",x"FF",x"D5",x"FF",x"D5",x"FF",x"D5",x"FF",x"D5",x"FF",x"D5",x"FF",x"D5",x"FF"),
		(x"D5",x"FF",x"D5",x"D5",x"D5",x"FF",x"D5",x"00",x"D5",x"FF",x"D5",x"D5",x"D5",x"FF",x"D5"),
		(x"FF",x"D5",x"FF",x"D5",x"FF",x"D5",x"FF",x"00",x"FF",x"D5",x"FF",x"D5",x"FF",x"D5",x"FF"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"FF",x"D5",x"FF",x"00",x"FF",x"D5",x"FF",x"D5",x"FF",x"D5",x"FF",x"00",x"FF",x"D5",x"FF"),
		(x"D5",x"FF",x"D5",x"00",x"D5",x"FF",x"D5",x"D5",x"D5",x"FF",x"D5",x"00",x"D5",x"FF",x"D5"),
		(x"FF",x"D5",x"FF",x"00",x"FF",x"D5",x"FF",x"D5",x"FF",x"D5",x"FF",x"00",x"FF",x"D5",x"FF"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"FF",x"D5",x"FF",x"D5",x"FF",x"D5",x"FF",x"00",x"FF",x"D5",x"FF",x"D5",x"FF",x"D5",x"FF"),
		(x"D5",x"FF",x"D5",x"D5",x"D5",x"FF",x"D5",x"00",x"D5",x"FF",x"D5",x"D5",x"D5",x"FF",x"D5"),
		(x"FF",x"D5",x"FF",x"D5",x"FF",x"D5",x"FF",x"00",x"FF",x"D5",x"FF",x"D5",x"FF",x"D5",x"FF"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"FF",x"D5",x"FF",x"00",x"FF",x"D5",x"FF",x"D5",x"FF",x"D5",x"FF",x"00",x"FF",x"D5",x"FF"),
		(x"D5",x"FF",x"D5",x"00",x"D5",x"FF",x"D5",x"D5",x"D5",x"FF",x"D5",x"00",x"D5",x"FF",x"D5")
	
	);
	
	constant bloque_G : ROM :=
	(
	
		(x"D5",x"D5",x"D5",x"D5",x"D5",x"D5",x"D5",x"D5",x"D5",x"D5",x"D5",x"D5",x"D5",x"D5",x"D5"),
		(x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"00",x"55",x"55",x"55",x"55",x"55",x"55",x"55"),
		(x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"00",x"55",x"55",x"55",x"55",x"55",x"55",x"55"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"55",x"55",x"55",x"00",x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"00",x"55",x"55",x"55"),
		(x"55",x"55",x"55",x"00",x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"00",x"55",x"55",x"55"),
		(x"55",x"55",x"55",x"00",x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"00",x"55",x"55",x"55"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"00",x"55",x"55",x"55",x"55",x"55",x"55",x"55"),
		(x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"00",x"55",x"55",x"55",x"55",x"55",x"55",x"55"),
		(x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"00",x"55",x"55",x"55",x"55",x"55",x"55",x"55"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"55",x"55",x"55",x"00",x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"00",x"55",x"55",x"55"),
		(x"55",x"55",x"55",x"00",x"55",x"55",x"55",x"55",x"55",x"55",x"55",x"00",x"55",x"55",x"55")
	
	);
	
	constant bloque_B : ROM :=
	(
	
		(x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA",x"AA"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00")
	
	);
	
begin

	dat_R <= bloque_R( dir_y )( dir_x );
	dat_G <= bloque_G( dir_y )( dir_x );
	dat_B <= bloque_B( dir_y )( dir_x );

end comp;