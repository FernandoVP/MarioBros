library ieee;

use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity koopa_ROM is

	Port(
	
		dir_y : in integer;
		dir_x : in integer;
		
		dat_R : out std_logic_vector( 7 downto 0 );
		dat_G : out std_logic_vector( 7 downto 0 );
		dat_B : out std_logic_vector( 7 downto 0 )
		
	);

end koopa_ROM;

architecture comp of koopa_ROM is

	type arreglo is array( 0 to 37 ) of std_logic_vector( 0 to 7 );

	type ROM is array( 0 to 37 ) of arreglo;

	constant koopa_R : ROM :=
	(
	
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"01",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"01",x"FF",x"FE",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"01",x"01",x"01",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"01",x"02",x"01",x"01",x"FF",x"FF",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"01",x"FF",x"FF",x"01",x"02",x"01",x"01",x"01",x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"FF",x"00",x"FF",x"00",x"01",x"FF",x"FF",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"01",x"02",x"01",x"FF",x"01",x"01",x"01",x"01",x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"01",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"01",x"01",x"FF",x"FF",x"FF",x"01",x"01",x"01",x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"01",x"01",x"FF",x"FF",x"FF",x"01",x"FF",x"01",x"00",x"01",x"01",x"FF",x"FF",x"01",x"01",x"01",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"FE",x"FF",x"FF",x"FF",x"01",x"01",x"FF",x"FF",x"01",x"01",x"01",x"01",x"FF",x"FF",x"01",x"01",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"FF",x"00",x"01",x"00",x"01",x"FF",x"FF",x"01",x"01",x"01",x"01",x"01",x"FF",x"FF",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"01",x"FF",x"FF",x"FE",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"01",x"01",x"01",x"01",x"FF",x"FE",x"FF",x"01",x"01",x"FF",x"FF",x"FF",x"01",x"01",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"01",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"01",x"01",x"00",x"02",x"FF",x"FF",x"FF",x"00",x"01",x"01",x"01",x"01",x"01",x"01",x"02",x"01",x"FF",x"FF",x"02",x"FF",x"00",x"01",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"01",x"01",x"01",x"01",x"02",x"01",x"01",x"FF",x"FF",x"FF",x"01",x"01",x"01",x"00",x"01",x"02",x"01",x"01",x"00",x"01",x"02",x"00",x"01",x"FF",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"02",x"02",x"02",x"01",x"FF",x"FF",x"FF",x"01",x"01",x"01",x"01",x"00",x"01",x"FF",x"FF",x"FF",x"01",x"01",x"01",x"01",x"00",x"00",x"01",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"02",x"01",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"01",x"01",x"FF",x"FF",x"FE",x"01",x"01",x"01",x"FF",x"FF",x"FF",x"01",x"00",x"00",x"00"),
		(x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"01",x"00",x"01",x"00",x"00",x"00",x"00",x"01",x"01",x"FF",x"FF",x"FF",x"FF",x"FF",x"01",x"01",x"FF",x"FF",x"01",x"01",x"00",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"FF",x"FF",x"FF",x"00",x"00",x"FF",x"00",x"FF",x"FF",x"FE",x"FF",x"FF",x"01",x"01",x"01",x"01",x"01",x"02",x"01",x"FF",x"FF",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"00",x"FE",x"FF",x"FF",x"00",x"FF",x"FF",x"FE",x"01",x"FE",x"01",x"01",x"01",x"02",x"00",x"01",x"01",x"01",x"01",x"FF",x"00",x"01",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"01",x"01",x"FF",x"01",x"01",x"02",x"FF",x"FF",x"FF",x"01",x"01",x"01",x"FF",x"FF",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FE",x"FF",x"01",x"01",x"FF",x"FF",x"01",x"01",x"FF",x"FF",x"FF",x"01",x"01",x"01",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"01",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"01",x"01",x"00",x"FF",x"FE",x"00",x"01",x"01",x"FF",x"FF",x"01",x"01",x"FF",x"FF",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"01",x"01",x"01",x"FF",x"FE",x"01",x"01",x"00",x"01",x"01",x"01",x"01",x"FF",x"FE",x"FF",x"01",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"01",x"01",x"00",x"01",x"01",x"FF",x"00",x"00",x"01",x"01",x"FE",x"FF",x"01",x"FF",x"FF",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"01",x"01",x"01",x"01",x"FF",x"FF",x"01",x"01",x"01",x"FF",x"00",x"01",x"FF",x"01",x"00",x"01",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"02",x"01",x"00",x"00",x"FF",x"FF",x"FF",x"00",x"01",x"00",x"01",x"00",x"01",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"02",x"01",x"01",x"01",x"01",x"FF",x"FF",x"FF",x"FF",x"01",x"01",x"01",x"01",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"FF",x"00",x"01",x"02",x"01",x"01",x"01",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"01",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00")
	
	);
	
	constant koopa_G : ROM :=
	(
	
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"02",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"01",x"00",x"A8",x"A8",x"FF",x"FF",x"FF",x"A0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"A8",x"A8",x"A8",x"FF",x"FF",x"A0",x"A0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"A8",x"A9",x"A8",x"A8",x"A0",x"A0",x"A8",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"A0",x"00",x"00",x"A8",x"FF",x"FF",x"A8",x"A9",x"A8",x"A8",x"A8",x"A8",x"A8",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"A0",x"00",x"A0",x"A7",x"A8",x"FF",x"FF",x"A8",x"A8",x"A9",x"A8",x"A9",x"A8",x"A8",x"A8",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"A0",x"A0",x"A0",x"FF",x"FF",x"FF",x"A8",x"A8",x"A8",x"A0",x"A8",x"A8",x"A8",x"A8",x"A9",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"01",x"00",x"00",x"9E",x"A0",x"9F",x"A0",x"FF",x"A7",x"A8",x"A8",x"A0",x"A0",x"9F",x"A8",x"A9",x"A8",x"A8",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"FF",x"FF",x"A0",x"A0",x"A8",x"A9",x"A0",x"A0",x"FF",x"A8",x"A0",x"A8",x"A9",x"A8",x"A8",x"FF",x"FF",x"A9",x"A8",x"A8",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"01",x"00",x"00",x"00",x"FF",x"00",x"A1",x"9F",x"A0",x"A0",x"A8",x"A8",x"A0",x"A0",x"A8",x"A8",x"A8",x"A8",x"FE",x"FF",x"A8",x"A8",x"FE",x"FF",x"A0",x"A9",x"00",x"01",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"FF",x"00",x"A8",x"00",x"A9",x"A0",x"A0",x"A9",x"A8",x"A8",x"A8",x"A8",x"FF",x"FF",x"A7",x"FF",x"FF",x"FF",x"A0",x"A0",x"A8",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"A0",x"A0",x"A0",x"A0",x"A0",x"A0",x"9F",x"A0",x"A0",x"A8",x"A8",x"A8",x"A8",x"FF",x"FE",x"FF",x"A8",x"A8",x"FF",x"A0",x"A0",x"A8",x"A8",x"FF",x"FF",x"A0",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"01",x"00",x"00",x"01",x"00",x"01",x"A0",x"A1",x"A0",x"A0",x"A0",x"A0",x"A0",x"A8",x"A8",x"A8",x"A8",x"FF",x"FF",x"FF",x"A7",x"A8",x"A8",x"A8",x"A8",x"A8",x"A8",x"A9",x"A9",x"A0",x"A0",x"A9",x"FF",x"00",x"00",x"00",x"00",x"01"),
		(x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"A8",x"A8",x"A8",x"A8",x"A8",x"A8",x"A8",x"A8",x"FF",x"FF",x"FF",x"A8",x"A8",x"A8",x"A7",x"A8",x"A9",x"A8",x"A8",x"A7",x"A8",x"A8",x"A7",x"A8",x"FF",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"A9",x"A9",x"A9",x"A9",x"A8",x"FF",x"FF",x"FF",x"A8",x"A8",x"A7",x"A8",x"A9",x"A8",x"FF",x"FF",x"FF",x"A8",x"A8",x"A9",x"A8",x"AA",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"A8",x"A8",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"A8",x"A9",x"FF",x"FF",x"9F",x"A8",x"A8",x"A9",x"FF",x"FE",x"FF",x"00",x"00",x"00",x"00"),
		(x"01",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"A8",x"A8",x"A0",x"A0",x"A0",x"FF",x"FF",x"A8",x"A8",x"A0",x"A0",x"A8",x"A8",x"A9",x"FF",x"FF",x"9E",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"A0",x"A0",x"A0",x"00",x"00",x"FF",x"00",x"A0",x"9F",x"A1",x"FE",x"FF",x"A8",x"A8",x"A8",x"A8",x"A8",x"A8",x"A8",x"A0",x"A0",x"00",x"01",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"A0",x"A0",x"FF",x"00",x"9F",x"A0",x"9F",x"00",x"FF",x"A0",x"A0",x"A8",x"FF",x"A8",x"A8",x"A8",x"A9",x"A9",x"A8",x"A9",x"A8",x"A8",x"FF",x"01",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"A2",x"A0",x"00",x"00",x"A1",x"A0",x"A0",x"A0",x"01",x"00",x"A8",x"A8",x"FF",x"A8",x"A8",x"A9",x"FF",x"FF",x"FF",x"A8",x"A8",x"A8",x"A0",x"FF",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"A1",x"FF",x"00",x"A0",x"9F",x"A0",x"A0",x"A0",x"9F",x"FF",x"A9",x"A8",x"FF",x"FF",x"A8",x"A8",x"FF",x"FF",x"A0",x"A8",x"A8",x"A8",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"A0",x"00",x"00",x"A0",x"A0",x"A0",x"A0",x"A1",x"A7",x"A9",x"A8",x"A7",x"FF",x"FE",x"A8",x"A8",x"A8",x"A0",x"A0",x"A8",x"A8",x"FF",x"FF",x"01",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FE",x"00",x"A0",x"A0",x"A0",x"A0",x"A0",x"A9",x"A8",x"A8",x"A9",x"FF",x"FE",x"A8",x"A8",x"A7",x"A8",x"A8",x"A8",x"A8",x"FF",x"FE",x"FF",x"01",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"01",x"00",x"00",x"FF",x"A0",x"A0",x"A0",x"00",x"A8",x"A8",x"A9",x"A8",x"A8",x"FF",x"AA",x"A9",x"A8",x"A8",x"FF",x"FF",x"A8",x"9F",x"A0",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"A8",x"A8",x"A8",x"A8",x"A8",x"FF",x"FF",x"A8",x"A8",x"A8",x"A0",x"A7",x"A8",x"A0",x"A8",x"00",x"01",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"A8",x"A8",x"A8",x"A9",x"A9",x"FF",x"FF",x"FE",x"A9",x"A8",x"A7",x"A9",x"A9",x"A8",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"A9",x"A8",x"A8",x"A8",x"A8",x"FF",x"FF",x"FF",x"FF",x"A8",x"A9",x"A8",x"A8",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"A0",x"A9",x"A9",x"A9",x"A8",x"A8",x"A8",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"01",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"A0",x"9F",x"A7",x"A7",x"A0",x"A1",x"A0",x"A0",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"A0",x"9F",x"A0",x"A0",x"A0",x"A0",x"A0",x"A0",x"A0",x"A0",x"FF",x"FF",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"A0",x"A0",x"FF",x"FF",x"A0",x"A0",x"A0",x"A0",x"01",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"A0",x"FF",x"FF",x"FF",x"A0",x"A0",x"A0",x"A0",x"A0",x"00",x"00",x"00")
		
	);
	
	constant koopa_B : ROM :=
	(
	
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FD",x"FF",x"FF",x"42",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"02",x"02",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"44",x"44",x"00",x"00",x"00",x"00",x"00",x"00",x"02",x"00",x"00",x"00",x"00",x"01",x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"02",x"FF",x"FF",x"00",x"01",x"00",x"00",x"44",x"44",x"02",x"00",x"00",x"02",x"00",x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"44",x"00",x"00",x"00",x"FF",x"FF",x"00",x"01",x"00",x"00",x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"44",x"00",x"44",x"00",x"00",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"02",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"02",x"00",x"44",x"42",x"44",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"44",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"02",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"01",x"00",x"00",x"43",x"42",x"44",x"44",x"FF",x"00",x"00",x"00",x"44",x"44",x"44",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"02",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"FF",x"FF",x"44",x"44",x"00",x"00",x"44",x"44",x"FF",x"00",x"42",x"00",x"00",x"00",x"00",x"FF",x"FF",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"44",x"44",x"44",x"44",x"00",x"00",x"44",x"44",x"00",x"00",x"00",x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"44",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"FF",x"00",x"00",x"00",x"00",x"44",x"44",x"00",x"02",x"00",x"00",x"00",x"FF",x"FF",x"00",x"FF",x"FF",x"FF",x"44",x"44",x"00",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"00",x"00",x"00",x"00",x"FF",x"FE",x"FF",x"00",x"02",x"FF",x"44",x"44",x"00",x"00",x"FF",x"FF",x"44",x"00",x"00",x"00",x"00",x"02",x"00",x"00"),
		(x"00",x"00",x"00",x"01",x"00",x"00",x"42",x"45",x"44",x"44",x"44",x"44",x"44",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"00",x"00",x"02",x"00",x"00",x"00",x"00",x"01",x"00",x"42",x"44",x"01",x"FF",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"01",x"01",x"00",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FD",x"FF",x"FF",x"FF",x"00",x"00",x"FF",x"FD",x"43",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"00",x"02",x"00",x"00"),
		(x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"44",x"44",x"44",x"FF",x"FF",x"00",x"00",x"44",x"44",x"00",x"00",x"00",x"FF",x"FF",x"43",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"44",x"44",x"44",x"00",x"00",x"FF",x"00",x"44",x"44",x"42",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"44",x"44",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"44",x"42",x"FF",x"02",x"43",x"44",x"44",x"00",x"FF",x"44",x"46",x"00",x"FF",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"45",x"42",x"00",x"02",x"45",x"44",x"44",x"44",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"01",x"FF",x"FF",x"FD",x"00",x"00",x"00",x"44",x"FF",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"45",x"FF",x"00",x"44",x"46",x"44",x"44",x"42",x"43",x"FF",x"00",x"00",x"FF",x"FF",x"00",x"00",x"FF",x"FF",x"44",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"44",x"00",x"00",x"44",x"44",x"44",x"44",x"45",x"00",x"00",x"00",x"00",x"FF",x"FF",x"00",x"00",x"00",x"44",x"44",x"00",x"00",x"FF",x"FF",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"44",x"44",x"44",x"44",x"44",x"00",x"00",x"00",x"00",x"FF",x"FE",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FE",x"FF",x"01",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"03",x"00",x"00",x"00",x"FF",x"44",x"44",x"44",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"01",x"00",x"00",x"00",x"FF",x"FF",x"00",x"44",x"44",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"00",x"00",x"00",x"44",x"00",x"00",x"45",x"00",x"00",x"01",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"44",x"00",x"00",x"01",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FD",x"FF",x"FF",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"42",x"44",x"00",x"00",x"46",x"45",x"44",x"44",x"FF",x"FF",x"FF",x"FF",x"FF",x"02",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"42",x"FF",x"FF",x"00",x"02",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"44",x"42",x"FF",x"FF",x"44",x"44",x"44",x"44",x"00",x"00",x"00",x"00"),
		(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"02",x"00",x"FF",x"FF",x"FF",x"44",x"FF",x"FF",x"FF",x"44",x"44",x"44",x"44",x"44",x"00",x"00",x"00")
		
	);
	
begin

	dat_R <= koopa_R( dir_y )( dir_x );
	dat_G <= koopa_G( dir_y )( dir_x );
	dat_B <= koopa_B( dir_y )( dir_x );

end comp;