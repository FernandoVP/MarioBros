library ieee;

use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity titulo_ROM is

	Port(
	
		dir_y : in integer;
		dir_x : in integer;
		
		dat_R : out std_logic_vector( 7 downto 0 );
		dat_G : out std_logic_vector( 7 downto 0 );
		dat_B : out std_logic_vector( 7 downto 0 )
		
	);

end titulo_ROM;

architecture comp of titulo_ROM is

	type arreglo is array( 0 to 175 ) of std_logic_vector( 0 to 7 );

	type ROM is array( 0 to 87 ) of arreglo;
	
	constant titulo_R : ROM :=
	(
	
		(x"FF",x"FF",x"FA",x"FF",x"FC",x"FD",x"FF",x"FE",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FB",x"F7",x"F8",x"FF",x"FF",x"FC",x"FC",x"FF"),
		(x"FF",x"FF",x"F7",x"FF",x"FF",x"FD",x"FF",x"F6",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FD",x"FF",x"FF",x"FF",x"FF",x"FB",x"FE",x"FF",x"FF"),
		(x"F6",x"FE",x"95",x"A1",x"9C",x"99",x"A3",x"9A",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"95",x"A4",x"94",x"8E",x"9B",x"98",x"90",x"99"),
		(x"F9",x"FF",x"A5",x"9F",x"91",x"91",x"86",x"9D",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"A1",x"9B",x"8F",x"9A",x"9A",x"9E",x"9B",x"A7"),
		(x"FF",x"FF",x"98",x"97",x"FF",x"FF",x"9F",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9E",x"91",x"9A",x"98",x"FF",x"FF",x"9E",x"8D"),
		(x"FF",x"F9",x"93",x"90",x"FF",x"FF",x"00",x"A0",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"A0",x"95",x"9E",x"A8",x"FF",x"E5",x"14",x"9A"),
		(x"FF",x"FF",x"A9",x"87",x"9E",x"00",x"02",x"9A",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"99",x"8F",x"8F",x"9C",x"95",x"04",x"00",x"9A"),
		(x"FD",x"F8",x"9C",x"99",x"9C",x"A3",x"99",x"93",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"A1",x"98",x"9A",x"A4",x"94",x"9D",x"9F",x"8D"),
		(x"FF",x"FD",x"9C",x"98",x"9A",x"98",x"9B",x"98",x"98",x"94",x"9E",x"9A",x"99",x"94",x"96",x"95",x"93",x"9D",x"97",x"9C",x"98",x"9B",x"9E",x"A1",x"A6",x"A0",x"94",x"99",x"99",x"99",x"A4",x"99",x"9E",x"91",x"98",x"96",x"8C",x"95",x"94",x"9F",x"9E",x"91",x"98",x"96",x"8C",x"95",x"94",x"9F",x"93",x"9D",x"97",x"9C",x"98",x"9B",x"9E",x"A1",x"98",x"94",x"9E",x"9A",x"99",x"94",x"96",x"95",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"9E",x"91",x"98",x"96",x"8C",x"95",x"94",x"9F",x"93",x"9D",x"97",x"9C",x"98",x"9B",x"9E",x"A1",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A"),
		(x"FF",x"FD",x"9C",x"98",x"9A",x"98",x"9B",x"98",x"99",x"9E",x"9F",x"93",x"95",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"87",x"96",x"97",x"91",x"97",x"F5",x"FB",x"FF",x"FF",x"FF",x"FF",x"8F",x"A4",x"FF",x"FF",x"FA",x"FF",x"FF",x"FF",x"8F",x"A4",x"FF",x"FF",x"FA",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"87",x"96",x"97",x"99",x"9E",x"9F",x"93",x"95",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"8F",x"A4",x"FF",x"FF",x"FA",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"87",x"96",x"97",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A"),
		(x"FF",x"FD",x"9C",x"98",x"9A",x"98",x"9B",x"98",x"99",x"9F",x"96",x"98",x"FF",x"FB",x"F3",x"FF",x"EF",x"F4",x"FF",x"F4",x"FB",x"FF",x"8D",x"9D",x"9A",x"8F",x"FF",x"FC",x"FF",x"F3",x"FA",x"F1",x"9B",x"93",x"FF",x"FF",x"F7",x"FF",x"F7",x"FA",x"9B",x"93",x"FF",x"FF",x"F7",x"FF",x"F7",x"FA",x"EF",x"F4",x"FF",x"F4",x"FB",x"FF",x"8D",x"9D",x"99",x"9F",x"96",x"98",x"FF",x"FB",x"F3",x"FF",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"9B",x"93",x"FF",x"FF",x"F7",x"FF",x"F7",x"FA",x"EF",x"F4",x"FF",x"F4",x"FB",x"FF",x"8D",x"9D",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A"),
		(x"FF",x"FD",x"9C",x"98",x"9A",x"98",x"9B",x"98",x"9E",x"9B",x"A3",x"8F",x"FC",x"F2",x"FE",x"F9",x"FF",x"FB",x"FB",x"FF",x"FC",x"FF",x"91",x"98",x"A3",x"9C",x"FF",x"FF",x"FF",x"FC",x"FF",x"FA",x"A0",x"9A",x"FF",x"FF",x"FB",x"FF",x"F8",x"FB",x"A0",x"9A",x"FF",x"FF",x"FB",x"FF",x"F8",x"FB",x"FF",x"FB",x"FB",x"FF",x"FC",x"FF",x"91",x"98",x"9E",x"9B",x"A3",x"8F",x"FC",x"F2",x"FE",x"F9",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"A0",x"9A",x"FF",x"FF",x"FB",x"FF",x"F8",x"FB",x"FF",x"FB",x"FB",x"FF",x"FC",x"FF",x"91",x"98",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A"),
		(x"FF",x"FD",x"9C",x"98",x"9A",x"98",x"9B",x"98",x"96",x"95",x"9F",x"FF",x"FE",x"FB",x"F7",x"FF",x"FF",x"FF",x"FE",x"FA",x"FF",x"FE",x"FF",x"95",x"94",x"9C",x"F9",x"FF",x"FF",x"F6",x"FF",x"F8",x"85",x"A8",x"FB",x"F9",x"FF",x"FF",x"FF",x"FE",x"85",x"A8",x"FB",x"F9",x"FF",x"FF",x"FF",x"FE",x"FF",x"FF",x"FE",x"FA",x"FF",x"FE",x"FF",x"95",x"96",x"95",x"9F",x"FF",x"FE",x"FB",x"F7",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"85",x"A8",x"FB",x"F9",x"FF",x"FF",x"FF",x"FE",x"FF",x"FF",x"FE",x"FA",x"FF",x"FE",x"FF",x"95",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A"),
		(x"FF",x"FD",x"9C",x"98",x"9A",x"98",x"9B",x"98",x"9A",x"94",x"8F",x"FF",x"FF",x"FA",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F9",x"FF",x"FF",x"86",x"98",x"97",x"FD",x"F6",x"FF",x"F9",x"FF",x"FF",x"11",x"91",x"FA",x"FD",x"F8",x"FF",x"FD",x"FC",x"11",x"91",x"FA",x"FD",x"F8",x"FF",x"FD",x"FC",x"FF",x"FF",x"FF",x"FF",x"F9",x"FF",x"FF",x"86",x"9A",x"94",x"8F",x"FF",x"FF",x"FA",x"FF",x"FF",x"FB",x"FB",x"FB",x"FB",x"FB",x"FB",x"FB",x"FB",x"11",x"91",x"FA",x"FD",x"F8",x"FF",x"FD",x"FC",x"FF",x"FF",x"FF",x"FF",x"F9",x"FF",x"FF",x"86",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A"),
		(x"FF",x"FD",x"9C",x"98",x"9A",x"98",x"9B",x"98",x"9F",x"96",x"FF",x"FF",x"FF",x"FF",x"FF",x"FB",x"FA",x"FB",x"FF",x"FF",x"F9",x"F5",x"FE",x"FF",x"9F",x"97",x"FF",x"FB",x"FF",x"FF",x"FF",x"FD",x"03",x"9A",x"FA",x"F7",x"F7",x"FD",x"FF",x"FD",x"03",x"9A",x"FA",x"F7",x"F7",x"FD",x"FF",x"FD",x"FA",x"FB",x"FF",x"FF",x"F9",x"F5",x"FE",x"FF",x"9F",x"96",x"FF",x"FF",x"FF",x"FF",x"FF",x"FB",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"03",x"9A",x"FA",x"F7",x"F7",x"FD",x"FF",x"FD",x"FA",x"FB",x"FF",x"FF",x"F9",x"F5",x"FE",x"FF",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A"),
		(x"FF",x"FD",x"9C",x"98",x"9A",x"98",x"9B",x"98",x"A0",x"91",x"FF",x"F7",x"FF",x"FF",x"F9",x"F9",x"F9",x"FF",x"FE",x"FF",x"FF",x"FF",x"FB",x"FF",x"9D",x"9B",x"FC",x"FF",x"FB",x"F5",x"FF",x"FA",x"00",x"9A",x"FF",x"FF",x"FF",x"FA",x"FF",x"FF",x"00",x"9A",x"FF",x"FF",x"FF",x"FA",x"FF",x"FF",x"F9",x"FF",x"FE",x"FF",x"FF",x"FF",x"FB",x"FF",x"A0",x"91",x"FF",x"F7",x"FF",x"FF",x"F9",x"F9",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"FE",x"00",x"9A",x"FF",x"FF",x"FF",x"FA",x"FF",x"FF",x"F9",x"FF",x"FE",x"FF",x"FF",x"FF",x"FB",x"FF",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A"),
		(x"FF",x"FD",x"9C",x"98",x"9A",x"98",x"9B",x"98",x"A1",x"A0",x"FA",x"FD",x"F7",x"FF",x"F3",x"FF",x"FF",x"FF",x"FC",x"FD",x"FF",x"FF",x"FD",x"FF",x"AB",x"95",x"FF",x"FF",x"FB",x"FF",x"FD",x"F7",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"FF",x"F3",x"FF",x"FF",x"FF",x"FF",x"F7",x"F8",x"7D",x"B1",x"FD",x"FF",x"FD",x"FF",x"FF",x"FB",x"FC",x"FF",x"FA",x"FF",x"FF",x"F7",x"FF",x"FF",x"00",x"9D",x"FF",x"F9",x"FD",x"FF",x"F0",x"FF",x"FA",x"FF",x"FB",x"EF",x"FD",x"FC",x"FF",x"F9",x"7A",x"B5",x"98",x"9B",x"96",x"9F",x"92",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A"),
		(x"FF",x"FD",x"9C",x"98",x"9A",x"98",x"9B",x"98",x"9C",x"8C",x"FE",x"FF",x"FF",x"FF",x"FF",x"FC",x"F7",x"08",x"00",x"00",x"00",x"03",x"08",x"02",x"87",x"9B",x"FA",x"FF",x"FF",x"FE",x"FF",x"FC",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"0E",x"FF",x"F8",x"F6",x"FF",x"FF",x"FB",x"FC",x"1A",x"95",x"FF",x"F9",x"FA",x"FF",x"FF",x"F9",x"00",x"04",x"03",x"00",x"00",x"00",x"01",x"00",x"00",x"99",x"FF",x"F9",x"FF",x"FF",x"F2",x"FF",x"04",x"FF",x"F8",x"FF",x"FF",x"FF",x"FF",x"FB",x"18",x"99",x"9A",x"95",x"94",x"A4",x"96",x"97",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A"),
		(x"FF",x"FD",x"9C",x"98",x"9A",x"98",x"9B",x"98",x"9E",x"8E",x"FF",x"FC",x"FB",x"FC",x"FF",x"F9",x"FC",x"F4",x"0D",x"00",x"07",x"07",x"00",x"00",x"11",x"98",x"FF",x"F4",x"FF",x"FF",x"FB",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"00",x"FF",x"FF",x"FB",x"FF",x"F7",x"FF",x"FF",x"06",x"99",x"FC",x"F6",x"FC",x"FF",x"FF",x"FF",x"05",x"F7",x"FF",x"FF",x"FF",x"FE",x"FF",x"00",x"00",x"96",x"FF",x"FD",x"FF",x"FF",x"F6",x"FF",x"00",x"F1",x"FF",x"FF",x"FF",x"F6",x"FF",x"FF",x"04",x"9C",x"96",x"91",x"97",x"9F",x"95",x"9F",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A"),
		(x"FF",x"FD",x"9C",x"98",x"9A",x"98",x"9B",x"98",x"A0",x"98",x"91",x"FF",x"EE",x"FD",x"FC",x"F9",x"FF",x"FE",x"FF",x"FF",x"07",x"00",x"00",x"00",x"06",x"91",x"FF",x"F8",x"FD",x"FF",x"FF",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"00",x"FF",x"F9",x"FB",x"FF",x"FB",x"FF",x"F3",x"02",x"96",x"F5",x"FD",x"FF",x"FC",x"FF",x"FE",x"04",x"FF",x"FF",x"F7",x"F8",x"FA",x"F9",x"0F",x"08",x"97",x"FF",x"FF",x"FF",x"FF",x"FA",x"FF",x"00",x"FD",x"F6",x"FD",x"FF",x"FC",x"FF",x"F7",x"00",x"99",x"91",x"9B",x"A1",x"9C",x"92",x"9D",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A"),
		(x"FF",x"FD",x"9C",x"98",x"9A",x"98",x"9B",x"98",x"91",x"A2",x"99",x"F6",x"FF",x"F7",x"FF",x"FD",x"FF",x"FF",x"F5",x"EF",x"FF",x"FF",x"07",x"00",x"0B",x"9B",x"FF",x"F9",x"FD",x"FF",x"F8",x"FE",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"02",x"FF",x"FE",x"F2",x"FF",x"FC",x"FF",x"04",x"01",x"97",x"FE",x"FF",x"FF",x"FD",x"FF",x"F8",x"00",x"F2",x"FF",x"FF",x"FF",x"FF",x"FE",x"0B",x"1A",x"85",x"F8",x"FF",x"FF",x"FF",x"FB",x"FD",x"10",x"F8",x"FB",x"FB",x"F9",x"F7",x"EE",x"0F",x"00",x"9A",x"9A",x"A0",x"9C",x"9D",x"99",x"98",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A"),
		(x"FF",x"FD",x"9C",x"98",x"9A",x"98",x"9B",x"98",x"96",x"99",x"A2",x"01",x"F7",x"ED",x"FF",x"FF",x"FF",x"F7",x"FF",x"FF",x"F1",x"FF",x"FF",x"96",x"84",x"9F",x"FF",x"FF",x"FE",x"FF",x"FC",x"FD",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"0D",x"FE",x"F4",x"FF",x"FF",x"F6",x"FC",x"00",x"09",x"9E",x"FF",x"FF",x"FD",x"F9",x"FF",x"FA",x"0F",x"FD",x"F9",x"F9",x"FF",x"F6",x"FF",x"7E",x"86",x"A5",x"FC",x"FF",x"FF",x"FA",x"FA",x"FF",x"06",x"FD",x"FC",x"F8",x"FF",x"FB",x"0F",x"00",x"07",x"A1",x"9F",x"A0",x"96",x"99",x"9A",x"98",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A"),
		(x"FF",x"FD",x"9C",x"98",x"9A",x"98",x"9B",x"98",x"9A",x"A0",x"91",x"0A",x"00",x"0B",x"FF",x"FF",x"F2",x"FF",x"F7",x"FF",x"FB",x"FA",x"FF",x"9F",x"91",x"9E",x"FC",x"FF",x"FB",x"FF",x"FF",x"FE",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"08",x"F8",x"FE",x"FF",x"FF",x"F6",x"0A",x"00",x"02",x"93",x"FC",x"FF",x"FF",x"F9",x"FF",x"FC",x"00",x"FF",x"FF",x"FE",x"FE",x"FF",x"FF",x"08",x"93",x"94",x"F7",x"FF",x"FF",x"FF",x"F9",x"FF",x"04",x"FF",x"FD",x"FF",x"FF",x"F3",x"F1",x"0B",x"00",x"95",x"98",x"9E",x"9C",x"9B",x"93",x"9C",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A"),
		(x"FF",x"FD",x"9C",x"98",x"9A",x"98",x"9B",x"98",x"8C",x"A6",x"98",x"95",x"00",x"14",x"00",x"00",x"FF",x"FD",x"FF",x"FF",x"FB",x"FC",x"FF",x"F7",x"A5",x"98",x"F6",x"FF",x"FA",x"FB",x"FF",x"F8",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"05",x"F6",x"FF",x"FF",x"FF",x"EC",x"00",x"0B",x"00",x"96",x"FF",x"F9",x"FB",x"F7",x"FF",x"FF",x"00",x"FF",x"FF",x"F8",x"F6",x"FF",x"FD",x"00",x"A5",x"99",x"FE",x"FF",x"F6",x"FF",x"FE",x"FF",x"00",x"F7",x"FE",x"FF",x"FA",x"F7",x"FF",x"FF",x"00",x"9A",x"9A",x"95",x"94",x"97",x"92",x"A5",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A"),
		(x"FF",x"FD",x"9C",x"98",x"9A",x"98",x"9B",x"98",x"9C",x"9D",x"8F",x"9F",x"07",x"00",x"0B",x"00",x"06",x"08",x"FB",x"FF",x"FF",x"FF",x"FE",x"F9",x"AA",x"98",x"FA",x"FA",x"FD",x"FC",x"FF",x"FF",x"0E",x"96",x"FC",x"FF",x"FF",x"FA",x"FF",x"F8",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"09",x"FB",x"FF",x"FF",x"FF",x"00",x"00",x"07",x"96",x"9F",x"FA",x"FF",x"FF",x"FD",x"FA",x"FF",x"11",x"78",x"0B",x"01",x"0A",x"00",x"00",x"01",x"A2",x"92",x"F7",x"FF",x"FF",x"FF",x"FF",x"F9",x"00",x"FF",x"F8",x"FA",x"FF",x"FE",x"FD",x"FF",x"A6",x"9A",x"99",x"9A",x"92",x"95",x"A0",x"9C",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A"),
		(x"FF",x"FD",x"9C",x"98",x"9A",x"98",x"9B",x"98",x"9E",x"96",x"FF",x"FF",x"F2",x"F7",x"FF",x"FF",x"ED",x"FA",x"FE",x"FC",x"FF",x"FF",x"F1",x"FF",x"99",x"98",x"F4",x"FF",x"FF",x"FB",x"FE",x"FC",x"EF",x"FF",x"FE",x"FE",x"FF",x"FF",x"FF",x"F9",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"00",x"8E",x"0B",x"00",x"01",x"00",x"00",x"14",x"9B",x"A2",x"F8",x"FF",x"FE",x"F5",x"FF",x"FF",x"FF",x"FF",x"FE",x"FA",x"FE",x"FE",x"F8",x"FF",x"9F",x"97",x"FF",x"FF",x"FC",x"FF",x"FF",x"F9",x"00",x"9A",x"FF",x"FC",x"FC",x"FD",x"FE",x"FF",x"92",x"94",x"93",x"A0",x"A1",x"95",x"9B",x"98",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A"),
		(x"FF",x"FD",x"9C",x"98",x"9A",x"98",x"9B",x"98",x"92",x"97",x"ED",x"FA",x"F4",x"FB",x"FF",x"FF",x"FF",x"FF",x"F7",x"FC",x"FE",x"FF",x"FF",x"FF",x"7F",x"A1",x"FF",x"FF",x"FC",x"FF",x"F8",x"FF",x"FF",x"F7",x"FF",x"FF",x"FF",x"FF",x"F5",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"0A",x"AC",x"00",x"04",x"0E",x"08",x"00",x"9B",x"90",x"94",x"FF",x"FD",x"FF",x"FB",x"FA",x"FE",x"FF",x"FB",x"FF",x"FC",x"FF",x"FE",x"FF",x"FF",x"A0",x"9A",x"FE",x"FF",x"FA",x"FF",x"FF",x"FC",x"06",x"88",x"FF",x"FF",x"FA",x"FF",x"FD",x"FE",x"85",x"A6",x"97",x"9B",x"9B",x"8E",x"9D",x"A1",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A"),
		(x"FF",x"FD",x"9C",x"98",x"9A",x"98",x"9B",x"98",x"97",x"9A",x"FF",x"F5",x"FB",x"FF",x"FE",x"FD",x"FF",x"FF",x"FD",x"FF",x"FF",x"F2",x"FF",x"F1",x"0E",x"98",x"FF",x"FF",x"FB",x"FD",x"FE",x"FF",x"FC",x"F6",x"FF",x"FF",x"F2",x"FF",x"F9",x"F9",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"00",x"98",x"00",x"0A",x"0A",x"0B",x"00",x"99",x"97",x"A3",x"FF",x"F8",x"FF",x"FB",x"FF",x"F5",x"F5",x"FF",x"F3",x"F7",x"FF",x"FC",x"FF",x"FE",x"93",x"9A",x"F9",x"FF",x"FC",x"FF",x"FC",x"FF",x"03",x"A3",x"F8",x"FF",x"F8",x"FF",x"FE",x"FD",x"1B",x"85",x"93",x"9C",x"A4",x"97",x"9E",x"97",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A"),
		(x"FF",x"FD",x"9C",x"98",x"9A",x"98",x"9B",x"98",x"A1",x"A8",x"A2",x"FF",x"FD",x"F3",x"FF",x"FA",x"FF",x"FF",x"F5",x"FF",x"FF",x"FA",x"F9",x"18",x"00",x"A0",x"8B",x"FF",x"FA",x"FF",x"FC",x"FF",x"FF",x"FF",x"FD",x"FF",x"F6",x"F8",x"FF",x"0A",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"00",x"A4",x"03",x"00",x"01",x"04",x"88",x"9D",x"94",x"9B",x"99",x"F7",x"FF",x"FF",x"FD",x"FF",x"FF",x"FE",x"FA",x"FF",x"FA",x"FF",x"FF",x"FF",x"81",x"AB",x"FF",x"FB",x"F7",x"FF",x"FB",x"FF",x"04",x"94",x"FF",x"FF",x"FF",x"FD",x"FF",x"FD",x"08",x"98",x"9F",x"9A",x"9E",x"94",x"9E",x"99",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A"),
		(x"FF",x"FD",x"9C",x"98",x"9A",x"98",x"9B",x"98",x"90",x"93",x"A6",x"FC",x"FC",x"FF",x"FF",x"F9",x"F1",x"FC",x"F5",x"FF",x"FF",x"F7",x"F5",x"06",x"00",x"9F",x"97",x"F4",x"FF",x"F7",x"FF",x"FF",x"F3",x"FF",x"FF",x"FD",x"FA",x"FF",x"F8",x"03",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"9A",x"8D",x"9C",x"98",x"93",x"A2",x"96",x"9B",x"9A",x"A1",x"E7",x"FF",x"FF",x"FF",x"FD",x"FF",x"F5",x"FF",x"FF",x"F4",x"F4",x"FA",x"F4",x"16",x"8C",x"FF",x"FD",x"FF",x"FF",x"FD",x"F8",x"06",x"99",x"FF",x"FF",x"FF",x"FB",x"FF",x"FC",x"00",x"97",x"9C",x"97",x"A1",x"94",x"98",x"9B",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A"),
		(x"FF",x"FD",x"9C",x"98",x"9A",x"98",x"9B",x"98",x"91",x"91",x"93",x"0A",x"F2",x"FF",x"F9",x"FB",x"FD",x"F7",x"FF",x"F9",x"FF",x"FD",x"0E",x"02",x"00",x"A2",x"90",x"0C",x"FF",x"F8",x"FF",x"FB",x"FF",x"FF",x"FF",x"F6",x"FE",x"FF",x"0D",x"00",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"16",x"86",x"9F",x"9E",x"9C",x"9A",x"A2",x"9E",x"99",x"9E",x"97",x"0D",x"FB",x"FF",x"FF",x"FA",x"FF",x"FF",x"FF",x"FF",x"FF",x"FD",x"FF",x"FB",x"07",x"9B",x"FF",x"F8",x"FB",x"FF",x"FE",x"FF",x"01",x"A0",x"F8",x"FB",x"FB",x"FD",x"FF",x"FE",x"00",x"98",x"9B",x"93",x"9F",x"95",x"95",x"9E",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A"),
		(x"FF",x"FD",x"9C",x"98",x"9A",x"98",x"9B",x"98",x"A4",x"A3",x"8B",x"02",x"FE",x"FF",x"FF",x"FF",x"FF",x"F6",x"FF",x"FA",x"F5",x"FD",x"04",x"00",x"02",x"96",x"A0",x"00",x"FF",x"F7",x"FF",x"F6",x"FA",x"FD",x"FF",x"F8",x"FF",x"FF",x"00",x"00",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"00",x"A0",x"96",x"99",x"9B",x"9D",x"9C",x"8F",x"9E",x"91",x"9B",x"04",x"FA",x"FC",x"FF",x"FA",x"FF",x"F6",x"FF",x"FF",x"F6",x"FF",x"FF",x"FC",x"00",x"97",x"FF",x"FD",x"FF",x"FF",x"F9",x"FC",x"05",x"90",x"FF",x"FF",x"FF",x"FF",x"FF",x"FA",x"00",x"9D",x"A2",x"93",x"9B",x"95",x"92",x"9F",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A"),
		(x"FF",x"FD",x"9C",x"98",x"9A",x"98",x"9B",x"98",x"8E",x"9C",x"A2",x"99",x"00",x"FF",x"FF",x"FF",x"FF",x"F3",x"F3",x"FF",x"FF",x"00",x"00",x"04",x"8E",x"9C",x"A2",x"99",x"00",x"FF",x"FF",x"FF",x"FF",x"F3",x"F3",x"FF",x"FF",x"00",x"00",x"04",x"90",x"98",x"FF",x"F7",x"F6",x"FD",x"FF",x"FF",x"00",x"9D",x"A2",x"93",x"9B",x"95",x"92",x"9F",x"8E",x"9C",x"A2",x"99",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"02",x"8E",x"FF",x"F5",x"FF",x"F8",x"F3",x"FF",x"02",x"8E",x"FF",x"F5",x"FF",x"F8",x"F3",x"FF",x"00",x"9D",x"A2",x"93",x"9B",x"95",x"92",x"9F",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A"),
		(x"FF",x"FD",x"9C",x"98",x"9A",x"98",x"9B",x"98",x"A1",x"9E",x"A7",x"8B",x"06",x"00",x"0C",x"00",x"05",x"00",x"08",x"10",x"00",x"00",x"00",x"04",x"A1",x"9E",x"A7",x"8B",x"06",x"00",x"0C",x"00",x"05",x"00",x"08",x"10",x"00",x"00",x"00",x"04",x"A1",x"A8",x"98",x"12",x"00",x"02",x"00",x"00",x"00",x"98",x"9B",x"93",x"9F",x"95",x"95",x"9E",x"A1",x"9E",x"A7",x"8B",x"06",x"00",x"0C",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"09",x"9A",x"94",x"0A",x"0D",x"09",x"00",x"03",x"09",x"9A",x"94",x"0A",x"0D",x"09",x"00",x"03",x"00",x"98",x"9B",x"93",x"9F",x"95",x"95",x"9E",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A"),
		(x"FF",x"FD",x"9C",x"98",x"9A",x"98",x"9B",x"98",x"9A",x"8C",x"9B",x"A7",x"A3",x"09",x"07",x"00",x"0A",x"0A",x"00",x"00",x"00",x"01",x"08",x"A3",x"9A",x"8C",x"9B",x"A7",x"A3",x"09",x"07",x"00",x"0A",x"0A",x"00",x"00",x"00",x"01",x"08",x"A3",x"9A",x"94",x"8F",x"02",x"00",x"06",x"04",x"00",x"00",x"97",x"9C",x"97",x"A1",x"94",x"98",x"9B",x"9A",x"8C",x"9B",x"A7",x"A3",x"09",x"07",x"00",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"96",x"9A",x"07",x"00",x"04",x"00",x"00",x"00",x"96",x"9A",x"07",x"00",x"04",x"00",x"00",x"00",x"97",x"9C",x"97",x"A1",x"94",x"98",x"9B",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A"),
		(x"FF",x"FD",x"9C",x"98",x"9A",x"98",x"9B",x"98",x"9E",x"92",x"9B",x"8D",x"95",x"03",x"01",x"01",x"0B",x"07",x"03",x"06",x"07",x"00",x"00",x"8A",x"9E",x"92",x"9B",x"8D",x"95",x"03",x"01",x"01",x"0B",x"07",x"03",x"06",x"07",x"00",x"00",x"8A",x"A3",x"8F",x"AC",x"00",x"01",x"0A",x"02",x"00",x"08",x"98",x"9F",x"9A",x"9E",x"94",x"9E",x"99",x"9E",x"92",x"9B",x"8D",x"95",x"03",x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"9A",x"94",x"09",x"00",x"01",x"00",x"02",x"00",x"9A",x"94",x"09",x"00",x"01",x"00",x"02",x"08",x"98",x"9F",x"9A",x"9E",x"94",x"9E",x"99",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A"),
		(x"FF",x"FD",x"9C",x"98",x"9A",x"98",x"9B",x"98",x"9F",x"9E",x"97",x"95",x"AA",x"90",x"07",x"00",x"00",x"00",x"00",x"03",x"00",x"08",x"92",x"9C",x"9F",x"9E",x"97",x"95",x"AA",x"90",x"07",x"00",x"00",x"00",x"00",x"03",x"00",x"08",x"92",x"9C",x"98",x"89",x"9A",x"00",x"04",x"07",x"00",x"00",x"1B",x"85",x"93",x"9C",x"A4",x"97",x"9E",x"97",x"9F",x"9E",x"97",x"95",x"AA",x"90",x"07",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"0B",x"9B",x"92",x"13",x"03",x"03",x"00",x"04",x"0B",x"9B",x"92",x"13",x"03",x"03",x"00",x"04",x"1B",x"85",x"93",x"9C",x"A4",x"97",x"9E",x"97",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A"),
		(x"FF",x"FD",x"9C",x"98",x"9A",x"98",x"9B",x"98",x"98",x"A2",x"A1",x"90",x"94",x"A4",x"94",x"9E",x"96",x"9C",x"9B",x"B0",x"98",x"98",x"A7",x"9E",x"98",x"A2",x"A1",x"90",x"94",x"A4",x"94",x"9E",x"96",x"9C",x"9B",x"B0",x"98",x"98",x"A7",x"9E",x"A2",x"96",x"AE",x"89",x"98",x"95",x"99",x"9E",x"85",x"A6",x"97",x"9B",x"9B",x"8E",x"9D",x"A1",x"98",x"A2",x"A1",x"90",x"94",x"A4",x"94",x"9E",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"9B",x"8D",x"9D",x"9F",x"94",x"9B",x"93",x"9B",x"AA",x"8D",x"9D",x"9F",x"94",x"9B",x"93",x"9B",x"AA",x"85",x"A6",x"97",x"9B",x"9B",x"8E",x"9D",x"A1",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A"),
		(x"FF",x"FD",x"9C",x"98",x"9A",x"98",x"9B",x"98",x"90",x"97",x"8A",x"8F",x"98",x"AA",x"90",x"93",x"9A",x"9A",x"8B",x"94",x"9B",x"91",x"90",x"97",x"90",x"97",x"8A",x"8F",x"98",x"AA",x"90",x"93",x"9A",x"9A",x"8B",x"94",x"9B",x"91",x"90",x"97",x"9F",x"90",x"9B",x"A3",x"98",x"96",x"9F",x"9C",x"92",x"94",x"93",x"A0",x"A1",x"95",x"9B",x"98",x"90",x"97",x"8A",x"8F",x"98",x"AA",x"90",x"93",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"93",x"9C",x"9D",x"95",x"A2",x"9E",x"99",x"99",x"93",x"9C",x"9D",x"95",x"A2",x"9E",x"99",x"99",x"92",x"94",x"93",x"A0",x"A1",x"95",x"9B",x"98",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A"),
		(x"FF",x"FD",x"9C",x"98",x"9A",x"98",x"9B",x"98",x"99",x"A5",x"97",x"A0",x"99",x"91",x"A2",x"9A",x"9A",x"9A",x"9F",x"91",x"9A",x"AE",x"97",x"99",x"99",x"A5",x"97",x"A0",x"99",x"91",x"A2",x"9A",x"9A",x"9A",x"9F",x"91",x"9A",x"AE",x"97",x"99",x"9D",x"92",x"98",x"9F",x"9F",x"93",x"8B",x"A3",x"A6",x"9A",x"99",x"9A",x"92",x"95",x"A0",x"9C",x"99",x"A5",x"97",x"A0",x"99",x"91",x"A2",x"9A",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"99",x"9E",x"9B",x"9B",x"90",x"9A",x"9B",x"96",x"96",x"9E",x"9B",x"9B",x"90",x"9A",x"9B",x"96",x"96",x"A6",x"9A",x"99",x"9A",x"92",x"95",x"A0",x"9C",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A"),
		(x"FF",x"FD",x"9C",x"98",x"9A",x"98",x"9B",x"98",x"98",x"94",x"9E",x"9A",x"99",x"94",x"96",x"95",x"8C",x"98",x"9B",x"98",x"9D",x"9A",x"92",x"9F",x"93",x"9D",x"97",x"9C",x"98",x"9B",x"9E",x"A1",x"98",x"94",x"9E",x"9A",x"99",x"94",x"96",x"95",x"93",x"9D",x"97",x"9C",x"98",x"9B",x"9E",x"A1",x"A6",x"A0",x"94",x"99",x"99",x"99",x"A4",x"99",x"93",x"9D",x"97",x"9C",x"98",x"9B",x"9E",x"A1",x"A6",x"A0",x"94",x"99",x"99",x"99",x"A4",x"99",x"9E",x"9C",x"9E",x"98",x"9C",x"9B",x"94",x"9B",x"93",x"9D",x"97",x"9C",x"98",x"9B",x"9E",x"A1",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"A6",x"A0",x"94",x"99",x"99",x"99",x"A4",x"99",x"93",x"9D",x"97",x"9C",x"98",x"9B",x"9E",x"A1",x"A6",x"A0",x"94",x"99",x"99",x"99",x"A4",x"99",x"93",x"9D",x"97",x"9C",x"98",x"9B",x"9E",x"A1",x"98",x"94",x"9E",x"9A",x"99",x"94",x"96",x"95",x"93",x"9D",x"97",x"9C",x"98",x"9B",x"9E",x"A1",x"98",x"94",x"9E",x"9A",x"99",x"94",x"96",x"95",x"93",x"9D",x"97",x"9C",x"98",x"9B",x"9E",x"A1",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A"),
		(x"FF",x"FD",x"9C",x"98",x"9A",x"98",x"9B",x"98",x"99",x"9E",x"9F",x"93",x"95",x"FF",x"FF",x"FF",x"FF",x"FF",x"8B",x"9B",x"A0",x"9B",x"9E",x"8E",x"FF",x"FF",x"FF",x"FF",x"FF",x"87",x"96",x"97",x"99",x"9E",x"9F",x"93",x"95",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"87",x"96",x"97",x"91",x"97",x"F5",x"FB",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"87",x"96",x"97",x"91",x"97",x"F5",x"FB",x"FF",x"FF",x"FF",x"FF",x"8A",x"99",x"9D",x"94",x"96",x"FF",x"FA",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"87",x"96",x"97",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"91",x"97",x"F5",x"FB",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"87",x"96",x"97",x"91",x"97",x"F5",x"FB",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"87",x"96",x"97",x"99",x"9E",x"9F",x"93",x"95",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"87",x"96",x"97",x"99",x"9E",x"9F",x"93",x"95",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"87",x"96",x"97",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A"),
		(x"FF",x"FD",x"9C",x"98",x"9A",x"98",x"9B",x"98",x"99",x"9F",x"96",x"98",x"FF",x"FB",x"F3",x"FF",x"FF",x"F5",x"FF",x"9A",x"8D",x"94",x"A0",x"FF",x"EF",x"F4",x"FF",x"F4",x"FB",x"FF",x"8D",x"9D",x"99",x"9F",x"96",x"98",x"FF",x"FB",x"F3",x"FF",x"EF",x"F4",x"FF",x"F4",x"FB",x"FF",x"8D",x"9D",x"9A",x"8F",x"FF",x"FC",x"FF",x"F3",x"FA",x"F1",x"EF",x"F4",x"FF",x"F4",x"FB",x"FF",x"8D",x"9D",x"9A",x"8F",x"FF",x"FC",x"FF",x"F3",x"FA",x"F1",x"9A",x"9D",x"9A",x"9A",x"FF",x"FF",x"F9",x"F2",x"EF",x"F4",x"FF",x"F4",x"FB",x"FF",x"8D",x"9D",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"8F",x"FF",x"FC",x"FF",x"F3",x"FA",x"F1",x"EF",x"F4",x"FF",x"F4",x"FB",x"FF",x"8D",x"9D",x"9A",x"8F",x"FF",x"FC",x"FF",x"F3",x"FA",x"F1",x"EF",x"F4",x"FF",x"F4",x"FB",x"FF",x"8D",x"9D",x"99",x"9F",x"96",x"98",x"FF",x"FB",x"F3",x"FF",x"EF",x"F4",x"FF",x"F4",x"FB",x"FF",x"8D",x"9D",x"99",x"9F",x"96",x"98",x"FF",x"FB",x"F3",x"FF",x"EF",x"F4",x"FF",x"F4",x"FB",x"FF",x"8D",x"9D",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A"),
		(x"FF",x"FD",x"9C",x"98",x"9A",x"98",x"9B",x"98",x"9E",x"9B",x"A3",x"8F",x"FC",x"F2",x"FE",x"F9",x"FF",x"F5",x"FF",x"8B",x"9D",x"A4",x"8F",x"FF",x"FF",x"FB",x"FB",x"FF",x"FC",x"FF",x"91",x"98",x"9E",x"9B",x"A3",x"8F",x"FC",x"F2",x"FE",x"F9",x"FF",x"FB",x"FB",x"FF",x"FC",x"FF",x"91",x"98",x"A3",x"9C",x"FF",x"FF",x"FF",x"FC",x"FF",x"FA",x"FF",x"FB",x"FB",x"FF",x"FC",x"FF",x"91",x"98",x"A3",x"9C",x"FF",x"FF",x"FF",x"FC",x"FF",x"FA",x"9D",x"9E",x"9D",x"8E",x"FF",x"F5",x"FF",x"FF",x"FF",x"FB",x"FB",x"FF",x"FC",x"FF",x"91",x"98",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"A3",x"9C",x"FF",x"FF",x"FF",x"FC",x"FF",x"FA",x"FF",x"FB",x"FB",x"FF",x"FC",x"FF",x"91",x"98",x"A3",x"9C",x"FF",x"FF",x"FF",x"FC",x"FF",x"FA",x"FF",x"FB",x"FB",x"FF",x"FC",x"FF",x"91",x"98",x"9E",x"9B",x"A3",x"8F",x"FC",x"F2",x"FE",x"F9",x"FF",x"FB",x"FB",x"FF",x"FC",x"FF",x"91",x"98",x"9E",x"9B",x"A3",x"8F",x"FC",x"F2",x"FE",x"F9",x"FF",x"FB",x"FB",x"FF",x"FC",x"FF",x"91",x"98",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A"),
		(x"FF",x"FD",x"9C",x"98",x"9A",x"98",x"9B",x"98",x"96",x"95",x"9F",x"FF",x"FE",x"FB",x"F7",x"FF",x"FA",x"FF",x"F8",x"FF",x"A0",x"99",x"FF",x"FF",x"FF",x"FF",x"FE",x"FA",x"FF",x"FE",x"FF",x"95",x"96",x"95",x"9F",x"FF",x"FE",x"FB",x"F7",x"FF",x"FF",x"FF",x"FE",x"FA",x"FF",x"FE",x"FF",x"95",x"94",x"9C",x"F9",x"FF",x"FF",x"F6",x"FF",x"F8",x"FF",x"FF",x"FE",x"FA",x"FF",x"FE",x"FF",x"95",x"94",x"9C",x"F9",x"FF",x"FF",x"F6",x"FF",x"F8",x"96",x"A3",x"9B",x"FF",x"F9",x"FD",x"FF",x"FF",x"FF",x"FF",x"FE",x"FA",x"FF",x"FE",x"FF",x"95",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"94",x"9C",x"F9",x"FF",x"FF",x"F6",x"FF",x"F8",x"FF",x"FF",x"FE",x"FA",x"FF",x"FE",x"FF",x"95",x"94",x"9C",x"F9",x"FF",x"FF",x"F6",x"FF",x"F8",x"FF",x"FF",x"FE",x"FA",x"FF",x"FE",x"FF",x"95",x"96",x"95",x"9F",x"FF",x"FE",x"FB",x"F7",x"FF",x"FF",x"FF",x"FE",x"FA",x"FF",x"FE",x"FF",x"95",x"96",x"95",x"9F",x"FF",x"FE",x"FB",x"F7",x"FF",x"FF",x"FF",x"FE",x"FA",x"FF",x"FE",x"FF",x"95",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A"),
		(x"FF",x"FD",x"9C",x"98",x"9A",x"98",x"9B",x"98",x"9A",x"94",x"8F",x"FF",x"FF",x"FA",x"FF",x"FF",x"FB",x"FF",x"FE",x"FF",x"9A",x"93",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F9",x"FF",x"FF",x"86",x"9A",x"94",x"8F",x"FF",x"FF",x"FA",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F9",x"FF",x"FF",x"86",x"98",x"97",x"FD",x"F6",x"FF",x"F9",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F9",x"FF",x"FF",x"86",x"98",x"97",x"FD",x"F6",x"FF",x"F9",x"FF",x"FF",x"0D",x"93",x"96",x"FF",x"FF",x"F6",x"FF",x"F6",x"FF",x"FF",x"FF",x"FF",x"F9",x"FF",x"FF",x"86",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"98",x"97",x"FD",x"F6",x"FF",x"F9",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F9",x"FF",x"FF",x"86",x"98",x"97",x"FD",x"F6",x"FF",x"F9",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F9",x"FF",x"FF",x"86",x"9A",x"94",x"8F",x"FF",x"FF",x"FA",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F9",x"FF",x"FF",x"86",x"9A",x"94",x"8F",x"FF",x"FF",x"FA",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F9",x"FF",x"FF",x"86",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A"),
		(x"FF",x"FD",x"9C",x"98",x"9A",x"98",x"9B",x"98",x"9F",x"96",x"FF",x"FF",x"FF",x"FF",x"FF",x"FB",x"FB",x"FF",x"FC",x"FF",x"FE",x"FF",x"FD",x"FF",x"FA",x"FB",x"FF",x"FF",x"F9",x"F5",x"FE",x"FF",x"9F",x"96",x"FF",x"FF",x"FF",x"FF",x"FF",x"FB",x"FA",x"FB",x"FF",x"FF",x"F9",x"F5",x"FE",x"FF",x"9F",x"97",x"FF",x"FB",x"FF",x"FF",x"FF",x"FD",x"FA",x"FB",x"FF",x"FF",x"F9",x"F5",x"FE",x"FF",x"9F",x"97",x"FF",x"FB",x"FF",x"FF",x"FF",x"FD",x"00",x"93",x"FF",x"FE",x"FF",x"F0",x"FF",x"F7",x"FA",x"FB",x"FF",x"FF",x"F9",x"F5",x"FE",x"FF",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9F",x"97",x"FF",x"FB",x"FF",x"FF",x"FF",x"FD",x"FA",x"FB",x"FF",x"FF",x"F9",x"F5",x"FE",x"FF",x"9F",x"97",x"FF",x"FB",x"FF",x"FF",x"FF",x"FD",x"FA",x"FB",x"FF",x"FF",x"F9",x"F5",x"FE",x"FF",x"9F",x"96",x"FF",x"FF",x"FF",x"FF",x"FF",x"FB",x"FA",x"FB",x"FF",x"FF",x"F9",x"F5",x"FE",x"FF",x"9F",x"96",x"FF",x"FF",x"FF",x"FF",x"FF",x"FB",x"FA",x"FB",x"FF",x"FF",x"F9",x"F5",x"FE",x"FF",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A"),
		(x"FF",x"FD",x"9C",x"98",x"9A",x"98",x"9B",x"98",x"A0",x"91",x"FF",x"F7",x"FF",x"FF",x"F9",x"F9",x"FF",x"F5",x"FF",x"FC",x"FC",x"FC",x"FF",x"F9",x"F9",x"FF",x"FE",x"FF",x"FF",x"FF",x"FB",x"FF",x"A0",x"91",x"FF",x"F7",x"FF",x"FF",x"F9",x"F9",x"F9",x"FF",x"FE",x"FF",x"FF",x"FF",x"FB",x"FF",x"9D",x"9B",x"FC",x"FF",x"FB",x"F5",x"FF",x"FA",x"F9",x"FF",x"FE",x"FF",x"FF",x"FF",x"FB",x"FF",x"9D",x"9B",x"FC",x"FF",x"FB",x"F5",x"FF",x"FA",x"00",x"A7",x"FF",x"F1",x"FF",x"FA",x"FD",x"FF",x"F9",x"FF",x"FE",x"FF",x"FF",x"FF",x"FB",x"FF",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9D",x"9B",x"FC",x"FF",x"FB",x"F5",x"FF",x"FA",x"F9",x"FF",x"FE",x"FF",x"FF",x"FF",x"FB",x"FF",x"9D",x"9B",x"FC",x"FF",x"FB",x"F5",x"FF",x"FA",x"F9",x"FF",x"FE",x"FF",x"FF",x"FF",x"FB",x"FF",x"A0",x"91",x"FF",x"F7",x"FF",x"FF",x"F9",x"F9",x"F9",x"FF",x"FE",x"FF",x"FF",x"FF",x"FB",x"FF",x"A0",x"91",x"FF",x"F7",x"FF",x"FF",x"F9",x"F9",x"F9",x"FF",x"FE",x"FF",x"FF",x"FF",x"FB",x"FF",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A"),
		(x"FF",x"FD",x"9C",x"98",x"9A",x"98",x"9B",x"98",x"9A",x"9D",x"FE",x"FA",x"FF",x"FD",x"FC",x"FF",x"F7",x"F4",x"FF",x"FB",x"FF",x"FC",x"FD",x"FF",x"F7",x"F4",x"FF",x"FB",x"FF",x"FC",x"FD",x"FF",x"7D",x"B1",x"FD",x"FF",x"FD",x"FF",x"FF",x"FB",x"F7",x"F4",x"FF",x"FB",x"FF",x"FC",x"FD",x"FF",x"7D",x"B1",x"FD",x"FF",x"FD",x"FF",x"FF",x"FB",x"F7",x"F4",x"FF",x"FB",x"FF",x"FC",x"FD",x"FF",x"7D",x"B1",x"FD",x"FF",x"FD",x"FF",x"FF",x"FB",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"F7",x"F4",x"FF",x"FB",x"FF",x"FC",x"FD",x"FF",x"7A",x"B5",x"98",x"9B",x"96",x"9F",x"92",x"9A",x"9A",x"9D",x"FE",x"FA",x"FF",x"FD",x"FC",x"FF",x"F7",x"F4",x"FF",x"FB",x"FF",x"FC",x"FD",x"FF",x"7D",x"B1",x"FD",x"FF",x"FD",x"FF",x"FF",x"FB",x"F7",x"F4",x"FF",x"FB",x"FF",x"FC",x"FD",x"FF",x"7D",x"B1",x"FD",x"FF",x"FD",x"FF",x"FF",x"FB",x"F7",x"F4",x"FF",x"FB",x"FF",x"FC",x"FD",x"FF",x"7D",x"B1",x"FD",x"FF",x"FD",x"FF",x"FF",x"FB",x"F7",x"F4",x"FF",x"FB",x"FF",x"FC",x"FD",x"FF",x"7A",x"B5",x"98",x"9B",x"96",x"9F",x"92",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A"),
		(x"FF",x"FD",x"9C",x"98",x"9A",x"98",x"9B",x"98",x"9A",x"9D",x"FE",x"FA",x"FF",x"FD",x"FC",x"FF",x"10",x"0A",x"FF",x"FC",x"FF",x"FB",x"FF",x"F7",x"10",x"0A",x"FF",x"FC",x"FF",x"FB",x"FF",x"F7",x"1A",x"95",x"FF",x"F9",x"FA",x"FF",x"FF",x"F9",x"10",x"0A",x"FF",x"FC",x"FF",x"FB",x"FF",x"F7",x"1A",x"95",x"FF",x"F9",x"FA",x"FF",x"FF",x"F9",x"10",x"0A",x"FF",x"FC",x"FF",x"FB",x"FF",x"F7",x"1A",x"95",x"FF",x"F9",x"FA",x"FF",x"FF",x"F9",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"10",x"0A",x"FF",x"FC",x"FF",x"FB",x"FF",x"F7",x"18",x"99",x"9A",x"95",x"94",x"A4",x"96",x"97",x"9A",x"9D",x"FE",x"FA",x"FF",x"FD",x"FC",x"FF",x"10",x"0A",x"FF",x"FC",x"FF",x"FB",x"FF",x"F7",x"1A",x"95",x"FF",x"F9",x"FA",x"FF",x"FF",x"F9",x"10",x"0A",x"FF",x"FC",x"FF",x"FB",x"FF",x"F7",x"1A",x"95",x"FF",x"F9",x"FA",x"FF",x"FF",x"F9",x"10",x"0A",x"FF",x"FC",x"FF",x"FB",x"FF",x"F7",x"1A",x"95",x"FF",x"F9",x"FA",x"FF",x"FF",x"F9",x"10",x"0A",x"FF",x"FC",x"FF",x"FB",x"FF",x"F7",x"18",x"99",x"9A",x"95",x"94",x"A4",x"96",x"97",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A"),
		(x"FF",x"FD",x"9C",x"98",x"9A",x"98",x"9B",x"98",x"9A",x"9D",x"FE",x"FA",x"FF",x"FD",x"FC",x"FF",x"01",x"00",x"FB",x"FF",x"F9",x"FD",x"FF",x"FF",x"01",x"00",x"FB",x"FF",x"F9",x"FD",x"FF",x"FF",x"06",x"99",x"FC",x"F6",x"FC",x"FF",x"FF",x"FF",x"01",x"00",x"FB",x"FF",x"F9",x"FD",x"FF",x"FF",x"06",x"99",x"FC",x"F6",x"FC",x"FF",x"FF",x"FF",x"01",x"00",x"FB",x"FF",x"F9",x"FD",x"FF",x"FF",x"06",x"99",x"FC",x"F6",x"FC",x"FF",x"FF",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"00",x"FB",x"FF",x"F9",x"FD",x"FF",x"FF",x"04",x"9C",x"96",x"91",x"97",x"9F",x"95",x"9F",x"9A",x"9D",x"FE",x"FA",x"FF",x"FD",x"FC",x"FF",x"01",x"00",x"FB",x"FF",x"F9",x"FD",x"FF",x"FF",x"06",x"99",x"FC",x"F6",x"FC",x"FF",x"FF",x"FF",x"01",x"00",x"FB",x"FF",x"F9",x"FD",x"FF",x"FF",x"06",x"99",x"FC",x"F6",x"FC",x"FF",x"FF",x"FF",x"01",x"00",x"FB",x"FF",x"F9",x"FD",x"FF",x"FF",x"06",x"99",x"FC",x"F6",x"FC",x"FF",x"FF",x"FF",x"01",x"00",x"FB",x"FF",x"F9",x"FD",x"FF",x"FF",x"04",x"9C",x"96",x"91",x"97",x"9F",x"95",x"9F",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A"),
		(x"FF",x"FD",x"9C",x"98",x"9A",x"98",x"9B",x"98",x"9A",x"9D",x"FE",x"FA",x"FF",x"FD",x"FC",x"FF",x"00",x"00",x"FF",x"FF",x"FA",x"FF",x"FF",x"FB",x"00",x"00",x"FF",x"FF",x"FA",x"FF",x"FF",x"FB",x"02",x"96",x"F5",x"FD",x"FF",x"FC",x"FF",x"FE",x"00",x"00",x"FF",x"FF",x"FA",x"FF",x"FF",x"FB",x"02",x"96",x"F5",x"FD",x"FF",x"FC",x"FF",x"FE",x"00",x"00",x"FF",x"FF",x"FA",x"FF",x"FF",x"FB",x"02",x"96",x"F5",x"FD",x"FF",x"FC",x"FF",x"FE",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"00",x"00",x"FF",x"FF",x"FA",x"FF",x"FF",x"FB",x"00",x"99",x"91",x"9B",x"A1",x"9C",x"92",x"9D",x"9A",x"9D",x"FE",x"FA",x"FF",x"FD",x"FC",x"FF",x"00",x"00",x"FF",x"FF",x"FA",x"FF",x"FF",x"FB",x"02",x"96",x"F5",x"FD",x"FF",x"FC",x"FF",x"FE",x"00",x"00",x"FF",x"FF",x"FA",x"FF",x"FF",x"FB",x"02",x"96",x"F5",x"FD",x"FF",x"FC",x"FF",x"FE",x"00",x"00",x"FF",x"FF",x"FA",x"FF",x"FF",x"FB",x"02",x"96",x"F5",x"FD",x"FF",x"FC",x"FF",x"FE",x"00",x"00",x"FF",x"FF",x"FA",x"FF",x"FF",x"FB",x"00",x"99",x"91",x"9B",x"A1",x"9C",x"92",x"9D",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A"),
		(x"FF",x"FD",x"9C",x"98",x"9A",x"98",x"9B",x"98",x"9A",x"9D",x"FE",x"FA",x"FF",x"FD",x"FC",x"FF",x"02",x"12",x"FF",x"FF",x"F6",x"FF",x"FF",x"F7",x"02",x"12",x"FF",x"FF",x"F6",x"FF",x"FF",x"F7",x"01",x"97",x"FE",x"FF",x"FF",x"FD",x"FF",x"F8",x"02",x"12",x"FF",x"FF",x"F6",x"FF",x"FF",x"F7",x"01",x"97",x"FE",x"FF",x"FF",x"FD",x"FF",x"F8",x"02",x"12",x"FF",x"FF",x"F6",x"FF",x"FF",x"F7",x"01",x"97",x"FE",x"FF",x"FF",x"FD",x"FF",x"F8",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"02",x"12",x"FF",x"FF",x"F6",x"FF",x"FF",x"F7",x"00",x"9A",x"9A",x"A0",x"9C",x"9D",x"99",x"98",x"9A",x"9D",x"FE",x"FA",x"FF",x"FD",x"FC",x"FF",x"02",x"12",x"FF",x"FF",x"F6",x"FF",x"FF",x"F7",x"01",x"97",x"FE",x"FF",x"FF",x"FD",x"FF",x"F8",x"02",x"12",x"FF",x"FF",x"F6",x"FF",x"FF",x"F7",x"01",x"97",x"FE",x"FF",x"FF",x"FD",x"FF",x"F8",x"02",x"12",x"FF",x"FF",x"F6",x"FF",x"FF",x"F7",x"01",x"97",x"FE",x"FF",x"FF",x"FD",x"FF",x"F8",x"02",x"12",x"FF",x"FF",x"F6",x"FF",x"FF",x"F7",x"00",x"9A",x"9A",x"A0",x"9C",x"9D",x"99",x"98",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A"),
		(x"FF",x"FD",x"9C",x"98",x"9A",x"98",x"9B",x"98",x"9A",x"9D",x"FE",x"FA",x"FF",x"FD",x"FC",x"FF",x"03",x"84",x"FD",x"FF",x"FD",x"FF",x"FD",x"FA",x"03",x"84",x"FD",x"FF",x"FD",x"FF",x"FD",x"FA",x"09",x"9E",x"FF",x"FF",x"FD",x"F9",x"FF",x"FA",x"03",x"84",x"FD",x"FF",x"FD",x"FF",x"FD",x"FA",x"09",x"9E",x"FF",x"FF",x"FD",x"F9",x"FF",x"FA",x"03",x"84",x"FD",x"FF",x"FD",x"FF",x"FD",x"FA",x"09",x"9E",x"FF",x"FF",x"FD",x"F9",x"FF",x"FA",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"03",x"84",x"FD",x"FF",x"FD",x"FF",x"FD",x"FA",x"07",x"A1",x"9F",x"A0",x"96",x"99",x"9A",x"98",x"9A",x"9D",x"FE",x"FA",x"FF",x"FD",x"FC",x"FF",x"03",x"84",x"FD",x"FF",x"FD",x"FF",x"FD",x"FA",x"09",x"9E",x"FF",x"FF",x"FD",x"F9",x"FF",x"FA",x"03",x"84",x"FD",x"FF",x"FD",x"FF",x"FD",x"FA",x"09",x"9E",x"FF",x"FF",x"FD",x"F9",x"FF",x"FA",x"03",x"84",x"FD",x"FF",x"FD",x"FF",x"FD",x"FA",x"09",x"9E",x"FF",x"FF",x"FD",x"F9",x"FF",x"FA",x"03",x"84",x"FD",x"FF",x"FD",x"FF",x"FD",x"FA",x"07",x"A1",x"9F",x"A0",x"96",x"99",x"9A",x"98",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A"),
		(x"FF",x"FD",x"9C",x"98",x"9A",x"98",x"9B",x"98",x"9A",x"9D",x"FE",x"FA",x"FF",x"FD",x"FC",x"FF",x"00",x"9F",x"FF",x"FF",x"F6",x"F8",x"FD",x"FF",x"00",x"9F",x"FF",x"FF",x"F6",x"F8",x"FD",x"FF",x"02",x"93",x"FC",x"FF",x"FF",x"F9",x"FF",x"FC",x"00",x"9F",x"FF",x"FF",x"F6",x"F8",x"FD",x"FF",x"02",x"93",x"FC",x"FF",x"FF",x"F9",x"FF",x"FC",x"00",x"9F",x"FF",x"FF",x"F6",x"F8",x"FD",x"FF",x"02",x"93",x"FC",x"FF",x"FF",x"F9",x"FF",x"FC",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"00",x"9F",x"FF",x"FF",x"F6",x"F8",x"FD",x"FF",x"00",x"95",x"98",x"9E",x"9C",x"9B",x"93",x"9C",x"9A",x"9D",x"FE",x"FA",x"FF",x"FD",x"FC",x"FF",x"00",x"9F",x"FF",x"FF",x"F6",x"F8",x"FD",x"FF",x"02",x"93",x"FC",x"FF",x"FF",x"F9",x"FF",x"FC",x"00",x"9F",x"FF",x"FF",x"F6",x"F8",x"FD",x"FF",x"02",x"93",x"FC",x"FF",x"FF",x"F9",x"FF",x"FC",x"00",x"9F",x"FF",x"FF",x"F6",x"F8",x"FD",x"FF",x"02",x"93",x"FC",x"FF",x"FF",x"F9",x"FF",x"FC",x"00",x"9F",x"FF",x"FF",x"F6",x"F8",x"FD",x"FF",x"00",x"95",x"98",x"9E",x"9C",x"9B",x"93",x"9C",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A"),
		(x"FF",x"FD",x"9C",x"98",x"9A",x"98",x"9B",x"98",x"9A",x"9D",x"FE",x"FA",x"FF",x"FD",x"FC",x"FF",x"00",x"9E",x"FB",x"FE",x"FF",x"FE",x"FF",x"FF",x"00",x"9E",x"FB",x"FE",x"FF",x"FE",x"FF",x"FF",x"00",x"96",x"FF",x"F9",x"FB",x"F7",x"FF",x"FF",x"00",x"9E",x"FB",x"FE",x"FF",x"FE",x"FF",x"FF",x"00",x"96",x"FF",x"F9",x"FB",x"F7",x"FF",x"FF",x"00",x"9E",x"FB",x"FE",x"FF",x"FE",x"FF",x"FF",x"00",x"96",x"FF",x"F9",x"FB",x"F7",x"FF",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"00",x"9E",x"FB",x"FE",x"FF",x"FE",x"FF",x"FF",x"00",x"9A",x"9A",x"95",x"94",x"97",x"92",x"A5",x"9A",x"9D",x"FE",x"FA",x"FF",x"FD",x"FC",x"FF",x"00",x"9E",x"FB",x"FE",x"FF",x"FE",x"FF",x"FF",x"00",x"96",x"FF",x"F9",x"FB",x"F7",x"FF",x"FF",x"00",x"9E",x"FB",x"FE",x"FF",x"FE",x"FF",x"FF",x"00",x"96",x"FF",x"F9",x"FB",x"F7",x"FF",x"FF",x"00",x"9E",x"FB",x"FE",x"FF",x"FE",x"FF",x"FF",x"00",x"96",x"FF",x"F9",x"FB",x"F7",x"FF",x"FF",x"00",x"9E",x"FB",x"FE",x"FF",x"FE",x"FF",x"FF",x"00",x"9A",x"9A",x"95",x"94",x"97",x"92",x"A5",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A"),
		(x"FF",x"FD",x"9C",x"98",x"9A",x"98",x"9B",x"98",x"9A",x"9D",x"FE",x"FA",x"FF",x"FD",x"FC",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"05",x"85",x"FF",x"FD",x"FE",x"F9",x"FF",x"F6",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"00",x"9A",x"98",x"9B",x"98",x"9A",x"95",x"9C",x"9A",x"9D",x"FE",x"FA",x"FF",x"FD",x"FC",x"FF",x"05",x"85",x"FF",x"FD",x"FE",x"F9",x"FF",x"F6",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"05",x"85",x"FF",x"FD",x"FE",x"F9",x"FF",x"F6",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"0A",x"9E",x"FE",x"F9",x"FD",x"FF",x"F1",x"FF",x"00",x"A5",x"F8",x"FB",x"FB",x"FF",x"EB",x"FF",x"00",x"9D",x"A2",x"93",x"9B",x"95",x"92",x"9F",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A"),
		(x"FF",x"FD",x"9C",x"98",x"9A",x"98",x"9B",x"98",x"9A",x"9D",x"FE",x"FA",x"FF",x"FD",x"FC",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"04",x"FF",x"FF",x"FC",x"FD",x"FF",x"FF",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"00",x"9A",x"98",x"9B",x"98",x"9A",x"95",x"9C",x"9A",x"9D",x"FE",x"FA",x"FF",x"FD",x"FC",x"FF",x"04",x"FF",x"FF",x"FC",x"FD",x"FF",x"FF",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"04",x"FF",x"FF",x"FC",x"FD",x"FF",x"FF",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"04",x"8A",x"FF",x"FD",x"FF",x"FE",x"FF",x"FD",x"FF",x"A2",x"90",x"04",x"09",x"00",x"07",x"04",x"00",x"98",x"9B",x"93",x"9F",x"95",x"95",x"9E",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A"),
		(x"FF",x"FD",x"9C",x"98",x"9A",x"98",x"9B",x"98",x"9A",x"9D",x"FE",x"FA",x"FF",x"FD",x"FC",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"0B",x"FE",x"FF",x"F2",x"FD",x"FD",x"FF",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"00",x"9A",x"98",x"9B",x"98",x"9A",x"95",x"9C",x"9A",x"9D",x"FE",x"FA",x"FF",x"FD",x"FC",x"FF",x"0B",x"FE",x"FF",x"F2",x"FD",x"FD",x"FF",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"0B",x"FE",x"FF",x"F2",x"FD",x"FD",x"FF",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"04",x"8C",x"FF",x"FA",x"FF",x"FA",x"FF",x"F9",x"FB",x"EB",x"9C",x"0D",x"06",x"05",x"0B",x"00",x"00",x"97",x"9C",x"97",x"A1",x"94",x"98",x"9B",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A"),
		(x"FF",x"FD",x"9C",x"98",x"9A",x"98",x"9B",x"98",x"9A",x"9D",x"FE",x"FA",x"FF",x"FD",x"FC",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"00",x"FF",x"FC",x"F7",x"FE",x"FD",x"FF",x"F2",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"00",x"9A",x"98",x"9B",x"98",x"9A",x"95",x"9C",x"9A",x"9D",x"FE",x"FA",x"FF",x"FD",x"FC",x"FF",x"00",x"FF",x"FC",x"F7",x"FE",x"FD",x"FF",x"F2",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"00",x"FF",x"FC",x"F7",x"FE",x"FD",x"FF",x"F2",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"07",x"96",x"96",x"FF",x"F3",x"FC",x"FB",x"FB",x"FF",x"FD",x"FF",x"EB",x"00",x"06",x"07",x"00",x"08",x"98",x"9F",x"9A",x"9E",x"94",x"9E",x"99",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A"),
		(x"FF",x"FD",x"9C",x"98",x"9A",x"98",x"9B",x"98",x"9A",x"9D",x"FE",x"FA",x"FF",x"FD",x"FC",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"F7",x"FF",x"FF",x"FE",x"F7",x"F2",x"06",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"00",x"9A",x"98",x"9B",x"98",x"9A",x"95",x"9C",x"9A",x"9D",x"FE",x"FA",x"FF",x"FD",x"FC",x"FF",x"01",x"F7",x"FF",x"FF",x"FE",x"F7",x"F2",x"06",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"F7",x"FF",x"FF",x"FE",x"F7",x"F2",x"06",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"00",x"A0",x"9E",x"F2",x"FF",x"F4",x"FF",x"FE",x"F4",x"FF",x"FF",x"FF",x"F2",x"F9",x"01",x"04",x"1B",x"85",x"93",x"9C",x"A4",x"97",x"9E",x"97",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A"),
		(x"FF",x"FD",x"9C",x"98",x"9A",x"98",x"9B",x"98",x"9A",x"9D",x"FE",x"FA",x"FF",x"FD",x"FC",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"00",x"FF",x"F9",x"FF",x"FF",x"FE",x"18",x"00",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"00",x"9A",x"98",x"9B",x"98",x"9A",x"95",x"9C",x"9A",x"9D",x"FE",x"FA",x"FF",x"FD",x"FC",x"FF",x"00",x"FF",x"F9",x"FF",x"FF",x"FE",x"18",x"00",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"00",x"FF",x"F9",x"FF",x"FF",x"FE",x"18",x"00",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"00",x"98",x"A6",x"00",x"FC",x"EA",x"FF",x"FF",x"FF",x"FF",x"F5",x"EF",x"F5",x"FF",x"F7",x"A1",x"85",x"A6",x"97",x"9B",x"9B",x"8E",x"9D",x"A1",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A"),
		(x"FF",x"FD",x"9C",x"98",x"9A",x"98",x"9B",x"98",x"9A",x"9D",x"FE",x"FA",x"FF",x"FD",x"FC",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"00",x"FF",x"FA",x"FF",x"FF",x"FC",x"F8",x"0A",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"00",x"9A",x"98",x"9B",x"98",x"9A",x"95",x"9C",x"9A",x"9D",x"FE",x"FA",x"FF",x"FD",x"FC",x"FF",x"00",x"FF",x"FA",x"FF",x"FF",x"FC",x"F8",x"0A",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"00",x"FF",x"FA",x"FF",x"FF",x"FC",x"F8",x"0A",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"00",x"9F",x"96",x"07",x"06",x"08",x"FF",x"FF",x"F8",x"FF",x"FF",x"F4",x"FF",x"FF",x"FC",x"8E",x"92",x"94",x"93",x"A0",x"A1",x"95",x"9B",x"98",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A"),
		(x"FF",x"FD",x"9C",x"98",x"9A",x"98",x"9B",x"98",x"9A",x"9D",x"FE",x"FA",x"FF",x"FD",x"FC",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"0C",x"FF",x"FA",x"F4",x"FF",x"FF",x"FF",x"F2",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"00",x"9A",x"98",x"9B",x"98",x"9A",x"95",x"9C",x"9A",x"9D",x"FE",x"FA",x"FF",x"FD",x"FC",x"FF",x"0C",x"FF",x"FA",x"F4",x"FF",x"FF",x"FF",x"F2",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"0C",x"FF",x"FA",x"F4",x"FF",x"FF",x"FF",x"F2",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"00",x"A5",x"9D",x"92",x"00",x"11",x"00",x"00",x"F5",x"FF",x"F2",x"FF",x"FF",x"F5",x"FF",x"FD",x"A6",x"9A",x"99",x"9A",x"92",x"95",x"A0",x"9C",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A"),
		(x"FF",x"FD",x"9C",x"98",x"9A",x"98",x"9B",x"98",x"9A",x"9D",x"FE",x"FA",x"FF",x"FD",x"FC",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"20",x"80",x"FC",x"FF",x"FE",x"FF",x"FC",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"00",x"FF",x"F8",x"FA",x"FF",x"FE",x"FD",x"FF",x"A5",x"99",x"FE",x"FF",x"F6",x"FF",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"00",x"9A",x"98",x"9B",x"98",x"9A",x"95",x"9C",x"9A",x"9D",x"FE",x"FA",x"FF",x"FD",x"FC",x"FF",x"08",x"F5",x"FF",x"F8",x"FF",x"FC",x"FD",x"FC",x"A5",x"99",x"FE",x"FF",x"F6",x"FF",x"FE",x"FF",x"00",x"FF",x"F8",x"FA",x"FF",x"FE",x"FD",x"FF",x"A5",x"99",x"FE",x"FF",x"F6",x"FF",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"03",x"AB",x"9B",x"8C",x"10",x"00",x"00",x"0C",x"06",x"00",x"FD",x"F9",x"FF",x"F3",x"FF",x"FE",x"A6",x"9A",x"99",x"9A",x"92",x"95",x"A0",x"9C",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A"),
		(x"FF",x"FD",x"9C",x"98",x"9A",x"98",x"9B",x"98",x"9A",x"9D",x"FE",x"FA",x"FF",x"FD",x"FC",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"FC",x"F3",x"FF",x"FC",x"FF",x"FF",x"FB",x"FE",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"00",x"9A",x"FF",x"FC",x"FC",x"FD",x"FE",x"FF",x"93",x"94",x"F7",x"FF",x"FF",x"FF",x"F9",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"00",x"9A",x"98",x"9B",x"98",x"9A",x"95",x"9C",x"9A",x"9D",x"FE",x"FA",x"FF",x"FD",x"FC",x"FF",x"00",x"0C",x"FF",x"FC",x"FF",x"F7",x"FF",x"FF",x"93",x"94",x"F7",x"FF",x"FF",x"FF",x"F9",x"FF",x"00",x"9A",x"FF",x"FC",x"FC",x"FD",x"FE",x"FF",x"93",x"94",x"F7",x"FF",x"FF",x"FF",x"F9",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"00",x"9A",x"FF",x"FF",x"F9",x"F0",x"FA",x"FD",x"00",x"11",x"FF",x"FF",x"FF",x"F4",x"F8",x"FF",x"92",x"94",x"93",x"A0",x"A1",x"95",x"9B",x"98",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A"),
		(x"FF",x"FD",x"9C",x"98",x"9A",x"98",x"9B",x"98",x"9A",x"9D",x"FE",x"FA",x"FF",x"FD",x"FC",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"FF",x"FB",x"FF",x"FF",x"FF",x"FF",x"FB",x"FE",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"06",x"88",x"FF",x"FF",x"FA",x"FF",x"FD",x"FE",x"86",x"A5",x"FC",x"FF",x"FF",x"FA",x"FA",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"00",x"9A",x"98",x"9B",x"98",x"9A",x"95",x"9C",x"9A",x"9D",x"FE",x"FA",x"FF",x"FD",x"FC",x"FF",x"00",x"00",x"FC",x"FB",x"FD",x"FF",x"FA",x"FF",x"86",x"A5",x"FC",x"FF",x"FF",x"FA",x"FA",x"FF",x"06",x"88",x"FF",x"FF",x"FA",x"FF",x"FD",x"FE",x"86",x"A5",x"FC",x"FF",x"FF",x"FA",x"FA",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"00",x"8A",x"FF",x"FB",x"FF",x"FF",x"FF",x"FD",x"07",x"0E",x"FA",x"FF",x"FF",x"F2",x"FE",x"FF",x"85",x"A6",x"97",x"9B",x"9B",x"8E",x"9D",x"A1",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A"),
		(x"FF",x"FD",x"9C",x"98",x"9A",x"98",x"9B",x"98",x"9A",x"9D",x"FE",x"FA",x"FF",x"FD",x"FC",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"F9",x"FF",x"FF",x"FF",x"F8",x"FC",x"FF",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"03",x"A3",x"F8",x"FF",x"F8",x"FF",x"FE",x"FD",x"1A",x"85",x"F8",x"FF",x"FF",x"FF",x"FB",x"FD",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"00",x"9A",x"98",x"9B",x"98",x"9A",x"95",x"9C",x"9A",x"9D",x"FE",x"FA",x"FF",x"FD",x"FC",x"FF",x"00",x"00",x"FF",x"FE",x"FF",x"FF",x"F4",x"FF",x"1A",x"85",x"F8",x"FF",x"FF",x"FF",x"FB",x"FD",x"03",x"A3",x"F8",x"FF",x"F8",x"FF",x"FE",x"FD",x"1A",x"85",x"F8",x"FF",x"FF",x"FF",x"FB",x"FD",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"10",x"A4",x"FB",x"FF",x"FF",x"FF",x"FC",x"F3",x"9B",x"00",x"FB",x"FF",x"FF",x"FF",x"F5",x"FF",x"1B",x"85",x"93",x"9C",x"A4",x"97",x"9E",x"97",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A"),
		(x"FF",x"FD",x"9C",x"98",x"9A",x"98",x"9B",x"98",x"9A",x"9D",x"FE",x"FA",x"FF",x"FD",x"FC",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"FB",x"FD",x"F6",x"FF",x"FF",x"FF",x"FC",x"FB",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"04",x"94",x"FF",x"FF",x"FF",x"FD",x"FF",x"FD",x"08",x"97",x"FF",x"FF",x"FF",x"FF",x"FA",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"00",x"9A",x"98",x"9B",x"98",x"9A",x"95",x"9C",x"9A",x"9D",x"FE",x"FA",x"FF",x"FD",x"FC",x"FF",x"07",x"0D",x"FE",x"FF",x"FF",x"FF",x"F8",x"FF",x"08",x"97",x"FF",x"FF",x"FF",x"FF",x"FA",x"FF",x"04",x"94",x"FF",x"FF",x"FF",x"FD",x"FF",x"FD",x"08",x"97",x"FF",x"FF",x"FF",x"FF",x"FA",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"00",x"98",x"F9",x"FF",x"FF",x"FB",x"FF",x"FB",x"92",x"06",x"F3",x"FF",x"EE",x"FF",x"FF",x"FF",x"08",x"98",x"9F",x"9A",x"9E",x"94",x"9E",x"99",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A"),
		(x"FF",x"FD",x"9C",x"98",x"9A",x"98",x"9B",x"98",x"9A",x"9D",x"FE",x"FA",x"FF",x"FD",x"FC",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"FF",x"FF",x"FA",x"FF",x"FC",x"FC",x"FC",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"06",x"99",x"FF",x"FF",x"FF",x"FB",x"FF",x"FC",x"00",x"96",x"FF",x"FD",x"FF",x"FF",x"F6",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"00",x"9A",x"98",x"9B",x"98",x"9A",x"95",x"9C",x"9A",x"9D",x"FE",x"FA",x"FF",x"FD",x"FC",x"FF",x"0A",x"82",x"FF",x"FF",x"FB",x"FF",x"FA",x"FD",x"00",x"96",x"FF",x"FD",x"FF",x"FF",x"F6",x"FF",x"06",x"99",x"FF",x"FF",x"FF",x"FB",x"FF",x"FC",x"00",x"96",x"FF",x"FD",x"FF",x"FF",x"F6",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"00",x"95",x"FC",x"FE",x"FC",x"F9",x"FF",x"FF",x"0A",x"8A",x"FF",x"FE",x"FF",x"FC",x"F9",x"FD",x"00",x"97",x"9C",x"97",x"A1",x"94",x"98",x"9B",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A"),
		(x"FF",x"FD",x"9C",x"98",x"9A",x"98",x"9B",x"98",x"9A",x"9D",x"FE",x"FA",x"FF",x"FD",x"FC",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"FC",x"FF",x"FD",x"FE",x"FE",x"FF",x"FD",x"F8",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"A0",x"F8",x"FB",x"FB",x"FD",x"FF",x"FE",x"00",x"99",x"FF",x"F9",x"FF",x"FF",x"F2",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"00",x"9A",x"98",x"9B",x"98",x"9A",x"95",x"9C",x"9A",x"9D",x"FE",x"FA",x"FF",x"FD",x"FC",x"FF",x"01",x"9D",x"FF",x"F8",x"FE",x"FF",x"FA",x"FF",x"00",x"99",x"FF",x"F9",x"FF",x"FF",x"F2",x"FF",x"01",x"A0",x"F8",x"FB",x"FB",x"FD",x"FF",x"FE",x"00",x"99",x"FF",x"F9",x"FF",x"FF",x"F2",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"03",x"9C",x"FF",x"FF",x"FA",x"FB",x"F9",x"FE",x"00",x"9D",x"FF",x"FF",x"FA",x"FD",x"FF",x"FE",x"00",x"98",x"9B",x"93",x"9F",x"95",x"95",x"9E",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A"),
		(x"FF",x"FD",x"9C",x"98",x"9A",x"98",x"9B",x"98",x"9A",x"9D",x"FE",x"FA",x"FF",x"FD",x"FC",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"FF",x"FF",x"FF",x"FD",x"FB",x"FE",x"FC",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"05",x"90",x"FF",x"FF",x"FF",x"FF",x"FF",x"FA",x"00",x"9D",x"FF",x"F9",x"FD",x"FF",x"F0",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"00",x"9A",x"98",x"9B",x"98",x"9A",x"95",x"9C",x"9A",x"9D",x"FE",x"FA",x"FF",x"FD",x"FC",x"FF",x"00",x"A9",x"F1",x"F6",x"F9",x"FF",x"FF",x"FC",x"00",x"9D",x"FF",x"F9",x"FD",x"FF",x"F0",x"FF",x"05",x"90",x"FF",x"FF",x"FF",x"FF",x"FF",x"FA",x"00",x"9D",x"FF",x"F9",x"FD",x"FF",x"F0",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"04",x"9D",x"FC",x"FE",x"FF",x"F8",x"FF",x"FC",x"0A",x"9D",x"F6",x"FF",x"FA",x"FC",x"FF",x"FF",x"00",x"9D",x"A2",x"93",x"9B",x"95",x"92",x"9F",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A"),
		(x"FF",x"FD",x"9C",x"98",x"9A",x"98",x"9B",x"98",x"9A",x"9D",x"FE",x"FA",x"FF",x"FD",x"FC",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"F7",x"F4",x"FF",x"FB",x"FF",x"FC",x"FD",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"A2",x"F8",x"FF",x"FE",x"FE",x"F7",x"FF",x"0E",x"96",x"FC",x"FF",x"FF",x"FA",x"FF",x"F8",x"00",x"9A",x"98",x"9B",x"98",x"9A",x"95",x"9C",x"9A",x"9D",x"FE",x"FA",x"FF",x"FD",x"FC",x"FF",x"00",x"91",x"FE",x"FD",x"FE",x"FF",x"FC",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"A2",x"F8",x"FF",x"FE",x"FE",x"F7",x"FF",x"0E",x"96",x"FC",x"FF",x"FF",x"FA",x"FF",x"F8",x"01",x"A2",x"F8",x"FF",x"FE",x"FE",x"F7",x"FF",x"0E",x"96",x"FC",x"FF",x"FF",x"FA",x"FF",x"F8",x"0A",x"A1",x"94",x"9A",x"99",x"99",x"9F",x"9B",x"9F",x"93",x"94",x"9D",x"9B",x"9C",x"9F",x"97"),
		(x"FF",x"FD",x"9C",x"98",x"9A",x"98",x"9B",x"98",x"9A",x"9D",x"FE",x"FA",x"FF",x"FD",x"FC",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"10",x"0A",x"FF",x"FC",x"FF",x"FB",x"FF",x"F7",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"02",x"A5",x"F8",x"FF",x"FC",x"F6",x"FD",x"FF",x"EF",x"FF",x"FE",x"FE",x"FF",x"FF",x"FF",x"F9",x"00",x"9A",x"98",x"9B",x"98",x"9A",x"95",x"9C",x"9A",x"9D",x"FE",x"FA",x"FF",x"FD",x"FC",x"FF",x"06",x"FF",x"FD",x"FA",x"FF",x"FF",x"FA",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"02",x"A5",x"F8",x"FF",x"FC",x"F6",x"FD",x"FF",x"EF",x"FF",x"FE",x"FE",x"FF",x"FF",x"FF",x"F9",x"02",x"A5",x"F8",x"FF",x"FC",x"F6",x"FD",x"FF",x"EF",x"FF",x"FE",x"FE",x"FF",x"FF",x"FF",x"F9",x"00",x"98",x"F4",x"FC",x"FF",x"FF",x"FF",x"FF",x"9E",x"97",x"9B",x"9D",x"98",x"9B",x"9E",x"99"),
		(x"FF",x"FD",x"9C",x"98",x"9A",x"98",x"9B",x"98",x"9A",x"9D",x"FE",x"FA",x"FF",x"FD",x"FC",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"00",x"FB",x"FF",x"F9",x"FD",x"FF",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"00",x"95",x"FF",x"FE",x"FF",x"FD",x"F7",x"FF",x"FF",x"F7",x"FF",x"FF",x"FF",x"FF",x"F5",x"FF",x"00",x"9A",x"98",x"9B",x"98",x"9A",x"95",x"9C",x"9A",x"9D",x"FE",x"FA",x"FF",x"FD",x"FC",x"FF",x"00",x"FF",x"FE",x"FF",x"F5",x"FF",x"FF",x"F7",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"00",x"95",x"FF",x"FE",x"FF",x"FD",x"F7",x"FF",x"FF",x"F7",x"FF",x"FF",x"FF",x"FF",x"F5",x"FF",x"00",x"95",x"FF",x"FE",x"FF",x"FD",x"F7",x"FF",x"FF",x"F7",x"FF",x"FF",x"FF",x"FF",x"F5",x"FF",x"01",x"8E",x"FF",x"FF",x"FF",x"F4",x"F5",x"F3",x"9F",x"9A",x"9B",x"99",x"98",x"9B",x"9B",x"9B"),
		(x"FF",x"FD",x"9C",x"98",x"9A",x"98",x"9B",x"98",x"9A",x"9D",x"FE",x"FA",x"FF",x"FD",x"FC",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"00",x"00",x"FF",x"FF",x"FA",x"FF",x"FF",x"FB",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"00",x"A4",x"FF",x"F7",x"FF",x"FC",x"FE",x"F7",x"FC",x"F6",x"FF",x"FF",x"F2",x"FF",x"F9",x"F9",x"00",x"9A",x"98",x"9B",x"98",x"9A",x"95",x"9C",x"9A",x"9D",x"FE",x"FA",x"FF",x"FD",x"FC",x"FF",x"02",x"FF",x"FA",x"FF",x"F5",x"FF",x"FF",x"EF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"00",x"A4",x"FF",x"F7",x"FF",x"FC",x"FE",x"F7",x"FC",x"F6",x"FF",x"FF",x"F2",x"FF",x"F9",x"F9",x"00",x"A4",x"FF",x"F7",x"FF",x"FC",x"FE",x"F7",x"FC",x"F6",x"FF",x"FF",x"F2",x"FF",x"F9",x"F9",x"08",x"9B",x"FF",x"FF",x"FF",x"FD",x"FF",x"FD",x"93",x"9A",x"96",x"96",x"99",x"9C",x"95",x"9E"),
		(x"FF",x"FD",x"9C",x"98",x"9A",x"98",x"9B",x"98",x"9A",x"9D",x"FE",x"FA",x"FF",x"FD",x"FC",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"02",x"12",x"FF",x"FF",x"F6",x"FF",x"FF",x"F7",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"00",x"9D",x"97",x"F7",x"FF",x"FF",x"FA",x"FF",x"FF",x"FF",x"FD",x"FF",x"F6",x"F8",x"FF",x"0A",x"00",x"9A",x"98",x"9B",x"98",x"9A",x"95",x"9C",x"9A",x"9D",x"FE",x"FA",x"FF",x"FD",x"FC",x"FF",x"02",x"F8",x"FE",x"FF",x"FD",x"FE",x"FE",x"0F",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"00",x"9D",x"97",x"F7",x"FF",x"FF",x"FA",x"FF",x"FF",x"FF",x"FD",x"FF",x"F6",x"F8",x"FF",x"0A",x"00",x"9D",x"97",x"F7",x"FF",x"FF",x"FA",x"FF",x"FF",x"FF",x"FD",x"FF",x"F6",x"F8",x"FF",x"0A",x"00",x"9D",x"F8",x"FF",x"FF",x"F8",x"FE",x"FA",x"80",x"AC",x"A3",x"94",x"94",x"9A",x"96",x"A0"),
		(x"FF",x"FD",x"9C",x"98",x"9A",x"98",x"9B",x"98",x"9A",x"9D",x"FE",x"FA",x"FF",x"FD",x"FC",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"03",x"84",x"FD",x"FF",x"FD",x"FF",x"FD",x"FA",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"9B",x"A0",x"E7",x"FF",x"FF",x"FE",x"FF",x"F3",x"FF",x"FF",x"FD",x"FA",x"FF",x"F8",x"03",x"00",x"9A",x"98",x"9B",x"98",x"9A",x"95",x"9C",x"9A",x"9D",x"FE",x"FA",x"FF",x"FD",x"FC",x"FF",x"00",x"FF",x"F9",x"FF",x"FB",x"FA",x"FB",x"03",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"9B",x"A0",x"E7",x"FF",x"FF",x"FE",x"FF",x"F3",x"FF",x"FF",x"FD",x"FA",x"FF",x"F8",x"03",x"01",x"9B",x"A0",x"E7",x"FF",x"FF",x"FE",x"FF",x"F3",x"FF",x"FF",x"FD",x"FA",x"FF",x"F8",x"03",x"00",x"97",x"FA",x"F7",x"FF",x"FB",x"FF",x"FF",x"15",x"8C",x"9F",x"95",x"9C",x"A1",x"96",x"96"),
		(x"FF",x"FD",x"9C",x"98",x"9A",x"98",x"9B",x"98",x"9A",x"9D",x"FE",x"FA",x"FF",x"FD",x"FC",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"00",x"9F",x"FF",x"FF",x"F6",x"F8",x"FD",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"03",x"A0",x"96",x"0D",x"FA",x"FF",x"FD",x"FC",x"FF",x"FF",x"FF",x"F6",x"FE",x"FF",x"0D",x"00",x"00",x"9A",x"98",x"9B",x"98",x"9A",x"95",x"9C",x"9A",x"9D",x"FE",x"FA",x"FF",x"FD",x"FC",x"FF",x"02",x"FF",x"F7",x"FE",x"FF",x"FF",x"0D",x"00",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"03",x"A0",x"96",x"0D",x"FA",x"FF",x"FD",x"FC",x"FF",x"FF",x"FF",x"F6",x"FE",x"FF",x"0D",x"00",x"03",x"A0",x"96",x"0D",x"FA",x"FF",x"FD",x"FC",x"FF",x"FF",x"FF",x"F6",x"FE",x"FF",x"0D",x"00",x"06",x"99",x"FF",x"FE",x"FF",x"FF",x"FF",x"FE",x"07",x"9C",x"A4",x"90",x"97",x"9C",x"98",x"9F"),
		(x"FF",x"FD",x"9C",x"98",x"9A",x"98",x"9B",x"98",x"9A",x"9D",x"FE",x"FA",x"FF",x"FD",x"FC",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"00",x"9E",x"FB",x"FE",x"FF",x"FE",x"FF",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"04",x"93",x"9A",x"05",x"F7",x"FD",x"FF",x"FC",x"FA",x"FD",x"FF",x"F8",x"FF",x"FF",x"00",x"00",x"00",x"9A",x"98",x"9B",x"98",x"9A",x"95",x"9C",x"9A",x"9D",x"FE",x"FA",x"FF",x"FD",x"FC",x"FF",x"00",x"FF",x"FE",x"FD",x"FF",x"FB",x"04",x"00",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"01",x"98",x"FE",x"FF",x"FE",x"FE",x"FE",x"FF",x"04",x"93",x"9A",x"05",x"F7",x"FD",x"FF",x"FC",x"FA",x"FD",x"FF",x"F8",x"FF",x"FF",x"00",x"00",x"04",x"93",x"9A",x"05",x"F7",x"FD",x"FF",x"FC",x"FA",x"FD",x"FF",x"F8",x"FF",x"FF",x"00",x"00",x"03",x"9A",x"FC",x"FF",x"FC",x"F5",x"FF",x"FC",x"00",x"98",x"9D",x"96",x"A5",x"9C",x"92",x"9B"),
		(x"FB",x"FF",x"95",x"A3",x"A1",x"9F",x"97",x"A2",x"90",x"98",x"FF",x"F7",x"F6",x"FD",x"FF",x"FF",x"02",x"8E",x"FF",x"F5",x"FF",x"F8",x"F3",x"FF",x"02",x"8E",x"FF",x"F5",x"FF",x"F8",x"F3",x"FF",x"02",x"8E",x"FF",x"F5",x"FF",x"F8",x"F3",x"FF",x"02",x"8E",x"FF",x"F5",x"FF",x"F8",x"F3",x"FF",x"02",x"8E",x"FF",x"F5",x"FF",x"F8",x"F3",x"FF",x"02",x"8E",x"FF",x"F5",x"FF",x"F8",x"F3",x"FF",x"02",x"8E",x"FF",x"F5",x"FF",x"F8",x"F3",x"FF",x"00",x"A3",x"96",x"A5",x"00",x"FF",x"FB",x"FF",x"FF",x"F3",x"F3",x"FF",x"FF",x"00",x"00",x"04",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"90",x"98",x"FF",x"F7",x"F6",x"FD",x"FF",x"FF",x"08",x"F7",x"FF",x"FF",x"FB",x"01",x"06",x"01",x"90",x"98",x"FF",x"F7",x"F6",x"FD",x"FF",x"FF",x"02",x"8E",x"FF",x"F5",x"FF",x"F8",x"F3",x"FF",x"00",x"A3",x"96",x"A5",x"00",x"FF",x"FB",x"FF",x"FF",x"F3",x"F3",x"FF",x"FF",x"00",x"00",x"04",x"8E",x"9C",x"A2",x"99",x"00",x"FF",x"FF",x"FF",x"FF",x"F3",x"F3",x"FF",x"FF",x"00",x"00",x"04",x"90",x"98",x"FF",x"F7",x"F6",x"FD",x"FF",x"FF",x"09",x"AB",x"8D",x"B0",x"9F",x"89",x"A4",x"94"),
		(x"FB",x"FF",x"A5",x"99",x"8F",x"97",x"92",x"97",x"A1",x"A8",x"98",x"12",x"00",x"02",x"00",x"00",x"09",x"9A",x"94",x"0A",x"0D",x"09",x"00",x"03",x"09",x"9A",x"94",x"0A",x"0D",x"09",x"00",x"03",x"09",x"9A",x"94",x"0A",x"0D",x"09",x"00",x"03",x"09",x"9A",x"94",x"0A",x"0D",x"09",x"00",x"03",x"09",x"9A",x"94",x"0A",x"0D",x"09",x"00",x"03",x"09",x"9A",x"94",x"0A",x"0D",x"09",x"00",x"03",x"09",x"9A",x"94",x"0A",x"0D",x"09",x"00",x"03",x"01",x"A0",x"84",x"90",x"03",x"00",x"04",x"00",x"05",x"00",x"08",x"10",x"00",x"00",x"00",x"04",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"A1",x"A8",x"98",x"12",x"00",x"02",x"00",x"00",x"00",x"A8",x"03",x"00",x"07",x"00",x"0F",x"00",x"A1",x"A8",x"98",x"12",x"00",x"02",x"00",x"00",x"09",x"9A",x"94",x"0A",x"0D",x"09",x"00",x"03",x"01",x"A0",x"84",x"90",x"03",x"00",x"04",x"00",x"05",x"00",x"08",x"10",x"00",x"00",x"00",x"04",x"A1",x"9E",x"A7",x"8B",x"06",x"00",x"0C",x"00",x"05",x"00",x"08",x"10",x"00",x"00",x"00",x"04",x"A1",x"A8",x"98",x"12",x"00",x"02",x"00",x"00",x"00",x"8D",x"9B",x"90",x"90",x"AD",x"9F",x"8B"),
		(x"F8",x"FF",x"94",x"8E",x"9C",x"9D",x"8E",x"9C",x"9A",x"94",x"8F",x"02",x"00",x"06",x"04",x"00",x"00",x"96",x"9A",x"07",x"00",x"04",x"00",x"00",x"00",x"96",x"9A",x"07",x"00",x"04",x"00",x"00",x"00",x"96",x"9A",x"07",x"00",x"04",x"00",x"00",x"00",x"96",x"9A",x"07",x"00",x"04",x"00",x"00",x"00",x"96",x"9A",x"07",x"00",x"04",x"00",x"00",x"00",x"96",x"9A",x"07",x"00",x"04",x"00",x"00",x"00",x"96",x"9A",x"07",x"00",x"04",x"00",x"00",x"00",x"A3",x"93",x"9E",x"98",x"01",x"07",x"00",x"0A",x"0A",x"00",x"00",x"00",x"01",x"08",x"A3",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"94",x"8F",x"02",x"00",x"06",x"04",x"00",x"08",x"97",x"00",x"08",x"03",x"04",x"08",x"9B",x"9A",x"94",x"8F",x"02",x"00",x"06",x"04",x"00",x"00",x"96",x"9A",x"07",x"00",x"04",x"00",x"00",x"00",x"A3",x"93",x"9E",x"98",x"01",x"07",x"00",x"0A",x"0A",x"00",x"00",x"00",x"01",x"08",x"A3",x"9A",x"8C",x"9B",x"A7",x"A3",x"09",x"07",x"00",x"0A",x"0A",x"00",x"00",x"00",x"01",x"08",x"A3",x"9A",x"94",x"8F",x"02",x"00",x"06",x"04",x"00",x"00",x"A1",x"98",x"99",x"8F",x"94",x"A5",x"9E"),
		(x"FF",x"FF",x"8D",x"99",x"9A",x"A3",x"96",x"AA",x"A3",x"8F",x"AC",x"00",x"01",x"0A",x"02",x"00",x"00",x"9A",x"94",x"09",x"00",x"01",x"00",x"02",x"00",x"9A",x"94",x"09",x"00",x"01",x"00",x"02",x"00",x"9A",x"94",x"09",x"00",x"01",x"00",x"02",x"00",x"9A",x"94",x"09",x"00",x"01",x"00",x"02",x"00",x"9A",x"94",x"09",x"00",x"01",x"00",x"02",x"00",x"9A",x"94",x"09",x"00",x"01",x"00",x"02",x"00",x"9A",x"94",x"09",x"00",x"01",x"00",x"02",x"07",x"9B",x"A5",x"9B",x"A6",x"08",x"02",x"00",x"0B",x"07",x"03",x"06",x"07",x"00",x"00",x"8A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"A3",x"8F",x"AC",x"00",x"01",x"0A",x"02",x"00",x"00",x"9B",x"0A",x"0D",x"00",x"01",x"00",x"94",x"A3",x"8F",x"AC",x"00",x"01",x"0A",x"02",x"00",x"00",x"9A",x"94",x"09",x"00",x"01",x"00",x"02",x"07",x"9B",x"A5",x"9B",x"A6",x"08",x"02",x"00",x"0B",x"07",x"03",x"06",x"07",x"00",x"00",x"8A",x"9E",x"92",x"9B",x"8D",x"95",x"03",x"01",x"01",x"0B",x"07",x"03",x"06",x"07",x"00",x"00",x"8A",x"A3",x"8F",x"AC",x"00",x"01",x"0A",x"02",x"00",x"07",x"9B",x"9B",x"93",x"8F",x"AC",x"9E",x"8E"),
		(x"FF",x"FE",x"9A",x"98",x"FF",x"FF",x"99",x"91",x"98",x"89",x"9A",x"00",x"04",x"07",x"00",x"00",x"0B",x"9B",x"92",x"13",x"03",x"03",x"00",x"04",x"0B",x"9B",x"92",x"13",x"03",x"03",x"00",x"04",x"0B",x"9B",x"92",x"13",x"03",x"03",x"00",x"04",x"0B",x"9B",x"92",x"13",x"03",x"03",x"00",x"04",x"0B",x"9B",x"92",x"13",x"03",x"03",x"00",x"04",x"0B",x"9B",x"92",x"13",x"03",x"03",x"00",x"04",x"0B",x"9B",x"92",x"13",x"03",x"03",x"00",x"04",x"06",x"8F",x"A3",x"9B",x"93",x"8A",x"07",x"03",x"00",x"00",x"00",x"03",x"00",x"08",x"92",x"9C",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"98",x"89",x"9A",x"00",x"04",x"07",x"00",x"00",x"00",x"AD",x"00",x"05",x"00",x"00",x"A0",x"9D",x"98",x"89",x"9A",x"00",x"04",x"07",x"00",x"00",x"0B",x"9B",x"92",x"13",x"03",x"03",x"00",x"04",x"06",x"8F",x"A3",x"9B",x"93",x"8A",x"07",x"03",x"00",x"00",x"00",x"03",x"00",x"08",x"92",x"9C",x"9F",x"9E",x"97",x"95",x"AA",x"90",x"07",x"00",x"00",x"00",x"00",x"03",x"00",x"08",x"92",x"9C",x"98",x"89",x"9A",x"00",x"04",x"07",x"00",x"00",x"00",x"A4",x"A8",x"99",x"FB",x"F3",x"A4",x"A4"),
		(x"FD",x"FA",x"98",x"A1",x"FF",x"E4",x"09",x"98",x"A2",x"96",x"AE",x"89",x"98",x"95",x"99",x"9E",x"8D",x"9D",x"9F",x"94",x"9B",x"93",x"9B",x"AA",x"8D",x"9D",x"9F",x"94",x"9B",x"93",x"9B",x"AA",x"8D",x"9D",x"9F",x"94",x"9B",x"93",x"9B",x"AA",x"8D",x"9D",x"9F",x"94",x"9B",x"93",x"9B",x"AA",x"8D",x"9D",x"9F",x"94",x"9B",x"93",x"9B",x"AA",x"8D",x"9D",x"9F",x"94",x"9B",x"93",x"9B",x"AA",x"8D",x"9D",x"9F",x"94",x"9B",x"93",x"9B",x"AA",x"84",x"96",x"97",x"8E",x"8F",x"A6",x"97",x"A8",x"96",x"9C",x"9B",x"B0",x"98",x"98",x"A7",x"9E",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"A2",x"96",x"AE",x"89",x"98",x"95",x"99",x"9E",x"92",x"9D",x"9B",x"97",x"92",x"93",x"9C",x"9B",x"A2",x"96",x"AE",x"89",x"98",x"95",x"99",x"9E",x"8D",x"9D",x"9F",x"94",x"9B",x"93",x"9B",x"AA",x"84",x"96",x"97",x"8E",x"8F",x"A6",x"97",x"A8",x"96",x"9C",x"9B",x"B0",x"98",x"98",x"A7",x"9E",x"98",x"A2",x"A1",x"90",x"94",x"A4",x"94",x"9E",x"96",x"9C",x"9B",x"B0",x"98",x"98",x"A7",x"9E",x"A2",x"96",x"AE",x"89",x"98",x"95",x"99",x"9E",x"8D",x"91",x"9C",x"9A",x"FE",x"F2",x"01",x"92"),
		(x"FE",x"FE",x"91",x"9F",x"9A",x"0E",x"00",x"A1",x"9F",x"90",x"9B",x"A3",x"98",x"96",x"9F",x"9C",x"93",x"9C",x"9D",x"95",x"A2",x"9E",x"99",x"99",x"93",x"9C",x"9D",x"95",x"A2",x"9E",x"99",x"99",x"93",x"9C",x"9D",x"95",x"A2",x"9E",x"99",x"99",x"93",x"9C",x"9D",x"95",x"A2",x"9E",x"99",x"99",x"93",x"9C",x"9D",x"95",x"A2",x"9E",x"99",x"99",x"93",x"9C",x"9D",x"95",x"A2",x"9E",x"99",x"99",x"93",x"9C",x"9D",x"95",x"A2",x"9E",x"99",x"99",x"A2",x"9F",x"A3",x"97",x"99",x"9B",x"8F",x"9D",x"9A",x"9A",x"8B",x"94",x"9B",x"91",x"90",x"97",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9F",x"90",x"9B",x"A3",x"98",x"96",x"9F",x"9C",x"98",x"9A",x"97",x"9A",x"A3",x"AC",x"A2",x"96",x"9F",x"90",x"9B",x"A3",x"98",x"96",x"9F",x"9C",x"93",x"9C",x"9D",x"95",x"A2",x"9E",x"99",x"99",x"A2",x"9F",x"A3",x"97",x"99",x"9B",x"8F",x"9D",x"9A",x"9A",x"8B",x"94",x"9B",x"91",x"90",x"97",x"90",x"97",x"8A",x"8F",x"98",x"AA",x"90",x"93",x"9A",x"9A",x"8B",x"94",x"9B",x"91",x"90",x"97",x"9F",x"90",x"9B",x"A3",x"98",x"96",x"9F",x"9C",x"A0",x"97",x"99",x"A9",x"8F",x"0F",x"03",x"95"),
		(x"FF",x"FF",x"97",x"A1",x"92",x"9E",x"97",x"8E",x"9D",x"92",x"98",x"9F",x"9F",x"93",x"8B",x"A3",x"9E",x"9B",x"9B",x"90",x"9A",x"9B",x"96",x"96",x"9E",x"9B",x"9B",x"90",x"9A",x"9B",x"96",x"96",x"9E",x"9B",x"9B",x"90",x"9A",x"9B",x"96",x"96",x"9E",x"9B",x"9B",x"90",x"9A",x"9B",x"96",x"96",x"9E",x"9B",x"9B",x"90",x"9A",x"9B",x"96",x"96",x"9E",x"9B",x"9B",x"90",x"9A",x"9B",x"96",x"96",x"9E",x"9B",x"9B",x"90",x"9A",x"9B",x"96",x"96",x"A2",x"97",x"8B",x"A3",x"A0",x"94",x"9E",x"9E",x"9A",x"9A",x"9F",x"91",x"9A",x"AE",x"97",x"99",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9A",x"9D",x"92",x"98",x"9F",x"9F",x"93",x"8B",x"A3",x"96",x"A6",x"9D",x"95",x"8E",x"99",x"95",x"93",x"9D",x"92",x"98",x"9F",x"9F",x"93",x"8B",x"A3",x"9E",x"9B",x"9B",x"90",x"9A",x"9B",x"96",x"96",x"A2",x"97",x"8B",x"A3",x"A0",x"94",x"9E",x"9E",x"9A",x"9A",x"9F",x"91",x"9A",x"AE",x"97",x"99",x"99",x"A5",x"97",x"A0",x"99",x"91",x"A2",x"9A",x"9A",x"9A",x"9F",x"91",x"9A",x"AE",x"97",x"99",x"9D",x"92",x"98",x"9F",x"9F",x"93",x"8B",x"A3",x"96",x"A5",x"8F",x"9D",x"99",x"9E",x"92",x"A5")
	
	);
	
	constant titulo_G : ROM :=
	(
		(x"01",x"00",x"04",x"0E",x"00",x"02",x"00",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"02",x"05",x"00",x"00",x"01",x"02",x"00",x"01"),
		(x"00",x"08",x"CF",x"C2",x"C7",x"CB",x"CE",x"CB",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"CD",x"D0",x"C2",x"CE",x"C4",x"CB",x"CB",x"C8",x"CF"),
		(x"00",x"D6",x"4D",x"50",x"52",x"54",x"49",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"4B",x"48",x"53",x"4E",x"54",x"4F",x"53",x"55",x"4C"),
		(x"08",x"C2",x"54",x"42",x"4B",x"4F",x"5B",x"4E",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4A",x"4B",x"54",x"5A",x"4B",x"4A",x"49",x"56"),
		(x"00",x"C6",x"4E",x"51",x"D4",x"C3",x"4F",x"50",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4D",x"53",x"4D",x"4A",x"CE",x"C4",x"51",x"4D"),
		(x"08",x"C7",x"4E",x"4E",x"C2",x"CB",x"00",x"47",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4F",x"4E",x"4A",x"50",x"4B",x"BF",x"D9",x"00",x"4B"),
		(x"00",x"D0",x"4F",x"5C",x"4E",x"00",x"02",x"4F",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"51",x"4D",x"58",x"51",x"50",x"00",x"06",x"4E"),
		(x"03",x"CD",x"4D",x"4A",x"52",x"4A",x"4E",x"53",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"4B",x"54",x"47",x"4D",x"4F",x"50",x"47",x"55"),
		(x"00",x"CD",x"4C",x"4F",x"4F",x"4F",x"4E",x"4F",x"4F",x"47",x"51",x"4F",x"51",x"4C",x"52",x"53",x"4C",x"54",x"4D",x"4C",x"4F",x"50",x"4D",x"4D",x"4B",x"4A",x"51",x"51",x"4C",x"4F",x"49",x"49",x"52",x"4C",x"54",x"4D",x"5B",x"53",x"51",x"48",x"52",x"4C",x"54",x"4D",x"5B",x"53",x"51",x"48",x"4C",x"54",x"4D",x"4C",x"4F",x"50",x"4D",x"4D",x"4F",x"47",x"51",x"4F",x"51",x"4C",x"52",x"53",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"50",x"52",x"4C",x"54",x"4D",x"5B",x"53",x"51",x"48",x"4C",x"54",x"4D",x"4C",x"4F",x"50",x"4D",x"4D",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E"),
		(x"00",x"CD",x"4C",x"4F",x"4F",x"4F",x"4E",x"4F",x"50",x"4C",x"4E",x"4B",x"55",x"C9",x"C9",x"C0",x"D2",x"C6",x"C6",x"CA",x"C6",x"50",x"54",x"4A",x"4E",x"58",x"C7",x"C8",x"D1",x"D0",x"C7",x"D0",x"48",x"60",x"C5",x"C9",x"CB",x"C1",x"C8",x"C9",x"48",x"60",x"C5",x"C9",x"CB",x"C1",x"C8",x"C9",x"D2",x"C6",x"C6",x"CA",x"C6",x"50",x"54",x"4A",x"50",x"4C",x"4E",x"4B",x"55",x"C9",x"C9",x"C0",x"CA",x"CA",x"CA",x"CA",x"CA",x"CA",x"CA",x"CA",x"48",x"60",x"C5",x"C9",x"CB",x"C1",x"C8",x"C9",x"D2",x"C6",x"C6",x"CA",x"C6",x"50",x"54",x"4A",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E"),
		(x"00",x"CD",x"4C",x"4F",x"4F",x"4F",x"4E",x"4F",x"4F",x"4F",x"40",x"53",x"C8",x"CE",x"C7",x"D2",x"C6",x"CE",x"D9",x"CA",x"CA",x"D0",x"50",x"54",x"53",x"4B",x"DB",x"CB",x"CD",x"CC",x"C9",x"D0",x"4F",x"49",x"CE",x"CB",x"D1",x"CE",x"D1",x"D1",x"4F",x"49",x"CE",x"CB",x"D1",x"CE",x"D1",x"D1",x"C6",x"CE",x"D9",x"CA",x"CA",x"D0",x"50",x"54",x"4F",x"4F",x"40",x"53",x"C8",x"CE",x"C7",x"D2",x"CE",x"CE",x"CE",x"CE",x"CE",x"CE",x"CE",x"CE",x"4F",x"49",x"CE",x"CB",x"D1",x"CE",x"D1",x"D1",x"C6",x"CE",x"D9",x"CA",x"CA",x"D0",x"50",x"54",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E"),
		(x"00",x"CD",x"4C",x"4F",x"4F",x"4F",x"4E",x"4F",x"54",x"48",x"4F",x"4F",x"CB",x"D4",x"D9",x"C8",x"D3",x"CB",x"CA",x"D4",x"CA",x"C8",x"4F",x"49",x"4A",x"48",x"C4",x"C7",x"C6",x"CC",x"D0",x"D1",x"52",x"43",x"CD",x"C8",x"CC",x"C7",x"C7",x"CD",x"52",x"43",x"CD",x"C8",x"CC",x"C7",x"C7",x"CD",x"D3",x"CB",x"CA",x"D4",x"CA",x"C8",x"4F",x"49",x"54",x"48",x"4F",x"4F",x"CB",x"D4",x"D9",x"C8",x"C8",x"C8",x"C8",x"C8",x"C8",x"C8",x"C8",x"C8",x"52",x"43",x"CD",x"C8",x"CC",x"C7",x"C7",x"CD",x"D3",x"CB",x"CA",x"D4",x"CA",x"C8",x"4F",x"49",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E"),
		(x"00",x"CD",x"4C",x"4F",x"4F",x"4F",x"4E",x"4F",x"52",x"47",x"57",x"C6",x"C9",x"D2",x"C9",x"CB",x"C7",x"CB",x"C4",x"C4",x"C9",x"C4",x"C6",x"50",x"47",x"56",x"C7",x"D1",x"CD",x"C9",x"C9",x"CB",x"52",x"57",x"CC",x"C8",x"CD",x"CF",x"C9",x"CC",x"52",x"57",x"CC",x"C8",x"CD",x"CF",x"C9",x"CC",x"C7",x"CB",x"C4",x"C4",x"C9",x"C4",x"C6",x"50",x"52",x"47",x"57",x"C6",x"C9",x"D2",x"C9",x"CB",x"CE",x"CE",x"CE",x"CE",x"CE",x"CE",x"CE",x"CE",x"52",x"57",x"CC",x"C8",x"CD",x"CF",x"C9",x"CC",x"C7",x"CB",x"C4",x"C4",x"C9",x"C4",x"C6",x"50",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E"),
		(x"00",x"CD",x"4C",x"4F",x"4F",x"4F",x"4E",x"4F",x"4F",x"4F",x"53",x"C4",x"C9",x"CB",x"CA",x"C6",x"CC",x"C6",x"D0",x"D1",x"CF",x"D4",x"C8",x"5B",x"52",x"57",x"D1",x"CA",x"D1",x"CE",x"C8",x"D2",x"00",x"46",x"D2",x"D1",x"CB",x"CA",x"C9",x"CC",x"00",x"46",x"D2",x"D1",x"CB",x"CA",x"C9",x"CC",x"CC",x"C6",x"D0",x"D1",x"CF",x"D4",x"C8",x"5B",x"4F",x"4F",x"53",x"C4",x"C9",x"CB",x"CA",x"C6",x"CB",x"CB",x"CB",x"CB",x"CB",x"CB",x"CB",x"CB",x"00",x"46",x"D2",x"D1",x"CB",x"CA",x"C9",x"CC",x"CC",x"C6",x"D0",x"D1",x"CF",x"D4",x"C8",x"5B",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E"),
		(x"00",x"CD",x"4C",x"4F",x"4F",x"4F",x"4E",x"4F",x"4E",x"54",x"CB",x"CA",x"CF",x"C9",x"D0",x"CD",x"CD",x"CC",x"CD",x"CC",x"CE",x"C7",x"CF",x"CB",x"4F",x"4C",x"CD",x"C6",x"CE",x"CD",x"C5",x"C9",x"03",x"4F",x"CE",x"C9",x"CB",x"D0",x"D0",x"CA",x"03",x"4F",x"CE",x"C9",x"CB",x"D0",x"D0",x"CA",x"CD",x"CC",x"CD",x"CC",x"CE",x"C7",x"CF",x"CB",x"4E",x"54",x"CB",x"CA",x"CF",x"C9",x"D0",x"CD",x"CB",x"CB",x"CB",x"CB",x"CB",x"CB",x"CB",x"CB",x"03",x"4F",x"CE",x"C9",x"CB",x"D0",x"D0",x"CA",x"CD",x"CC",x"CD",x"CC",x"CE",x"C7",x"CF",x"CB",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E"),
		(x"00",x"CD",x"4C",x"4F",x"4F",x"4F",x"4E",x"4F",x"47",x"52",x"CE",x"C7",x"CE",x"C8",x"C6",x"D2",x"CC",x"D2",x"C6",x"CB",x"CB",x"CE",x"C8",x"CB",x"4C",x"52",x"CA",x"CF",x"C9",x"CA",x"CE",x"CF",x"04",x"47",x"CC",x"C9",x"CB",x"C9",x"CA",x"CA",x"04",x"47",x"CC",x"C9",x"CB",x"C9",x"CA",x"CA",x"CC",x"D2",x"C6",x"CB",x"CB",x"CE",x"C8",x"CB",x"47",x"52",x"CE",x"C7",x"CE",x"C8",x"C6",x"D2",x"CB",x"CB",x"CB",x"CB",x"CB",x"CB",x"CB",x"CB",x"04",x"47",x"CC",x"C9",x"CB",x"C9",x"CA",x"CA",x"CC",x"D2",x"C6",x"CB",x"CB",x"CE",x"C8",x"CB",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E"),
		(x"00",x"CD",x"4C",x"4F",x"4F",x"4F",x"4E",x"4F",x"45",x"52",x"CC",x"CE",x"CD",x"C6",x"CD",x"CF",x"C8",x"CB",x"CC",x"CF",x"CF",x"CC",x"C9",x"C9",x"53",x"45",x"CF",x"C4",x"CB",x"CE",x"CB",x"CF",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"C7",x"CB",x"D2",x"CE",x"C8",x"CD",x"CB",x"D1",x"53",x"50",x"C6",x"CF",x"CC",x"CD",x"CA",x"CE",x"CA",x"CB",x"D1",x"C9",x"C8",x"CD",x"C7",x"CC",x"03",x"4F",x"C9",x"CE",x"CD",x"CE",x"D0",x"CA",x"CF",x"C5",x"D2",x"CC",x"CB",x"CD",x"CD",x"CD",x"53",x"4E",x"4A",x"52",x"4D",x"51",x"4D",x"51",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E"),
		(x"00",x"CD",x"4C",x"4F",x"4F",x"4F",x"4E",x"4F",x"53",x"57",x"C3",x"D0",x"D2",x"CC",x"C6",x"CB",x"D4",x"00",x"00",x"08",x"06",x"00",x"00",x"04",x"4C",x"53",x"CF",x"CC",x"D1",x"C6",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"CE",x"C8",x"C7",x"C9",x"D1",x"CD",x"C4",x"00",x"41",x"CF",x"CD",x"C9",x"CF",x"CC",x"C8",x"07",x"00",x"06",x"00",x"01",x"08",x"00",x"04",x"03",x"4D",x"C6",x"CC",x"CE",x"CD",x"CF",x"CA",x"00",x"D1",x"C4",x"CA",x"C7",x"CF",x"D2",x"CB",x"00",x"40",x"52",x"50",x"4B",x"53",x"4E",x"4C",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E"),
		(x"00",x"CD",x"4C",x"4F",x"4F",x"4F",x"4E",x"4F",x"4F",x"56",x"CA",x"C8",x"D3",x"CC",x"CA",x"CA",x"CB",x"C6",x"00",x"03",x"00",x"00",x"05",x"06",x"00",x"56",x"D3",x"C6",x"D3",x"C8",x"CA",x"CF",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"08",x"C5",x"D2",x"D3",x"C3",x"C9",x"CB",x"CB",x"00",x"51",x"D2",x"C9",x"C9",x"C8",x"C8",x"CE",x"04",x"C0",x"C3",x"CF",x"C5",x"C8",x"D6",x"00",x"01",x"50",x"CB",x"CC",x"CC",x"CA",x"D1",x"C8",x"08",x"C5",x"D5",x"C6",x"C3",x"C5",x"CA",x"CC",x"00",x"4F",x"56",x"4C",x"4B",x"4D",x"4B",x"52",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E"),
		(x"00",x"CD",x"4C",x"4F",x"4F",x"4F",x"4E",x"4F",x"4C",x"4A",x"51",x"CC",x"CA",x"CC",x"C7",x"D2",x"D1",x"CF",x"C5",x"CD",x"00",x"03",x"04",x"05",x"03",x"4D",x"CB",x"CD",x"CD",x"C5",x"CF",x"C9",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"06",x"C2",x"CF",x"D0",x"CB",x"CF",x"CB",x"CD",x"03",x"52",x"C8",x"CD",x"D2",x"C5",x"C7",x"CD",x"00",x"CF",x"CD",x"CA",x"CE",x"CD",x"C8",x"02",x"00",x"53",x"D3",x"CB",x"C8",x"C9",x"D3",x"C8",x"00",x"CC",x"C8",x"CC",x"CE",x"D5",x"CD",x"C4",x"03",x"50",x"4D",x"4F",x"54",x"49",x"4A",x"50",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E"),
		(x"00",x"CD",x"4C",x"4F",x"4F",x"4F",x"4E",x"4F",x"4C",x"51",x"4D",x"C5",x"D1",x"CC",x"CF",x"D0",x"C7",x"C8",x"D4",x"D1",x"C7",x"D9",x"00",x"01",x"00",x"4C",x"D1",x"C6",x"CC",x"CE",x"CC",x"CD",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"C4",x"D9",x"C1",x"C8",x"CD",x"C8",x"01",x"00",x"4D",x"CB",x"CC",x"CB",x"C8",x"D0",x"C8",x"03",x"CF",x"D1",x"C8",x"C7",x"CF",x"CB",x"00",x"00",x"40",x"CA",x"CB",x"CC",x"CC",x"CF",x"C6",x"03",x"C5",x"D5",x"D1",x"C4",x"D1",x"CD",x"00",x"00",x"4C",x"4E",x"4F",x"4D",x"4C",x"53",x"4C",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E"),
		(x"00",x"CD",x"4C",x"4F",x"4F",x"4F",x"4E",x"4F",x"52",x"4D",x"56",x"00",x"CD",x"D7",x"C1",x"BF",x"D3",x"C7",x"C7",x"C3",x"CA",x"CE",x"C2",x"4F",x"5D",x"4D",x"C4",x"CE",x"CB",x"C9",x"CD",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"CE",x"CD",x"D0",x"CA",x"C9",x"D3",x"05",x"04",x"51",x"CD",x"CA",x"C6",x"C8",x"D4",x"C9",x"00",x"CA",x"CC",x"CD",x"D3",x"C5",x"D5",x"5A",x"54",x"5C",x"D1",x"CA",x"C7",x"C6",x"CB",x"D1",x"00",x"CC",x"D1",x"C3",x"CB",x"D0",x"00",x"03",x"04",x"4F",x"51",x"4E",x"49",x"4C",x"56",x"4C",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E"),
		(x"00",x"CD",x"4C",x"4F",x"4F",x"4F",x"4E",x"4F",x"52",x"49",x"4F",x"00",x"01",x"00",x"D5",x"CE",x"CF",x"D5",x"C7",x"DC",x"CF",x"CA",x"C6",x"52",x"4C",x"4C",x"CA",x"C8",x"CE",x"CA",x"CB",x"CE",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"CC",x"CE",x"C9",x"C8",x"D1",x"00",x"01",x"01",x"47",x"C7",x"CD",x"D1",x"CC",x"CC",x"C8",x"03",x"CF",x"CC",x"CB",x"CC",x"C6",x"C2",x"00",x"4E",x"44",x"CC",x"CF",x"CE",x"CF",x"C9",x"C8",x"06",x"D0",x"CD",x"C7",x"CB",x"C8",x"D3",x"00",x"01",x"46",x"4B",x"50",x"53",x"4F",x"4E",x"4C",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E"),
		(x"00",x"CD",x"4C",x"4F",x"4F",x"4F",x"4E",x"4F",x"55",x"47",x"53",x"4E",x"0A",x"00",x"00",x"07",x"C9",x"C7",x"CB",x"C6",x"C9",x"CC",x"D4",x"C8",x"4F",x"4E",x"D1",x"CE",x"CE",x"C8",x"CF",x"C7",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"05",x"CA",x"C9",x"C9",x"CB",x"CE",x"09",x"00",x"02",x"51",x"CF",x"C9",x"CE",x"CA",x"C8",x"CD",x"02",x"C5",x"C7",x"CB",x"D1",x"CC",x"C6",x"07",x"54",x"46",x"D4",x"C8",x"C3",x"D0",x"CE",x"CB",x"02",x"C5",x"CC",x"D2",x"C7",x"D1",x"CD",x"C8",x"02",x"50",x"53",x"4D",x"4F",x"4E",x"4A",x"51",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E"),
		(x"00",x"CD",x"4C",x"4F",x"4F",x"4F",x"4E",x"4F",x"4A",x"50",x"50",x"4A",x"00",x"02",x"00",x"03",x"00",x"00",x"CA",x"CC",x"C8",x"C5",x"D6",x"C7",x"4B",x"4C",x"D2",x"D0",x"C5",x"D0",x"CF",x"CC",x"00",x"4A",x"CD",x"D1",x"C6",x"C7",x"C5",x"D2",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"D4",x"C2",x"CF",x"C8",x"02",x"06",x"01",x"4B",x"4B",x"CA",x"CD",x"C9",x"D3",x"C5",x"CB",x"00",x"60",x"00",x"00",x"06",x"00",x"03",x"01",x"4E",x"4C",x"D1",x"C8",x"CC",x"C8",x"CB",x"CC",x"00",x"CF",x"C8",x"C9",x"CE",x"CF",x"C8",x"CE",x"52",x"48",x"58",x"4A",x"47",x"54",x"4D",x"4F",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E"),
		(x"00",x"CD",x"4C",x"4F",x"4F",x"4F",x"4E",x"4F",x"52",x"48",x"D0",x"C7",x"D0",x"D2",x"CC",x"D4",x"CB",x"D7",x"CD",x"CB",x"CC",x"CA",x"C0",x"CF",x"4F",x"4B",x"C6",x"D1",x"CB",x"CB",x"CF",x"C3",x"CD",x"C7",x"CC",x"C9",x"C8",x"CF",x"CA",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"02",x"43",x"07",x"02",x"00",x"0C",x"05",x"00",x"54",x"52",x"C7",x"D1",x"C7",x"CB",x"CF",x"CC",x"C7",x"C9",x"C5",x"CC",x"C5",x"C8",x"CC",x"CD",x"4D",x"4D",x"D5",x"C8",x"CA",x"C9",x"CB",x"CD",x"00",x"55",x"CF",x"CA",x"CB",x"CE",x"C9",x"D0",x"4D",x"47",x"50",x"50",x"52",x"53",x"48",x"4C",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E"),
		(x"00",x"CD",x"4C",x"4F",x"4F",x"4F",x"4E",x"4F",x"51",x"55",x"C9",x"D2",x"CE",x"C6",x"C7",x"C6",x"CB",x"C8",x"C6",x"CB",x"CF",x"D3",x"CC",x"CF",x"55",x"52",x"CF",x"C2",x"C9",x"D1",x"CD",x"C9",x"D3",x"CE",x"CA",x"CB",x"D2",x"CA",x"C4",x"D0",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"01",x"4A",x"06",x"00",x"00",x"01",x"01",x"50",x"4D",x"47",x"CB",x"D0",x"CC",x"CF",x"CA",x"CF",x"D3",x"C3",x"D1",x"D2",x"CD",x"C9",x"D1",x"C6",x"53",x"4B",x"D0",x"CA",x"CD",x"CA",x"C9",x"CD",x"07",x"41",x"D1",x"D2",x"C8",x"D0",x"C7",x"CB",x"53",x"5E",x"53",x"4B",x"4B",x"4A",x"4C",x"54",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E"),
		(x"00",x"CD",x"4C",x"4F",x"4F",x"4F",x"4E",x"4F",x"4F",x"50",x"CD",x"CF",x"D5",x"D4",x"CC",x"CD",x"C2",x"CA",x"D0",x"CC",x"CC",x"CA",x"CA",x"C8",x"01",x"49",x"CA",x"C8",x"CB",x"C8",x"D4",x"C5",x"C3",x"CD",x"CD",x"CA",x"CA",x"D3",x"C4",x"D5",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"03",x"50",x"06",x"02",x"00",x"00",x"01",x"4D",x"54",x"57",x"C3",x"CD",x"CC",x"CB",x"D0",x"C9",x"C8",x"D8",x"C8",x"CC",x"CD",x"CB",x"D0",x"C5",x"52",x"48",x"C8",x"CA",x"D1",x"CC",x"C7",x"CF",x"00",x"58",x"C6",x"CF",x"C6",x"D1",x"C8",x"CC",x"00",x"42",x"4C",x"4C",x"51",x"50",x"50",x"4A",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E"),
		(x"00",x"CD",x"4C",x"4F",x"4F",x"4F",x"4E",x"4F",x"4B",x"52",x"49",x"C6",x"CD",x"BE",x"CB",x"CE",x"D5",x"C9",x"CA",x"C6",x"CB",x"D0",x"C9",x"00",x"04",x"52",x"4C",x"C9",x"C8",x"CE",x"D0",x"C7",x"D0",x"CD",x"C4",x"CF",x"D0",x"C5",x"CF",x"00",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"4C",x"0F",x"04",x"05",x"00",x"4F",x"55",x"4C",x"4E",x"4D",x"D3",x"C4",x"CC",x"C6",x"D3",x"CA",x"C4",x"C5",x"CE",x"C5",x"CD",x"C8",x"CF",x"51",x"5B",x"D1",x"CA",x"CC",x"CA",x"CB",x"D0",x"00",x"48",x"CA",x"CD",x"CB",x"CC",x"CB",x"CD",x"00",x"56",x"56",x"4C",x"4B",x"4D",x"52",x"4C",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E"),
		(x"00",x"CD",x"4C",x"4F",x"4F",x"4F",x"4E",x"4F",x"4C",x"4C",x"4D",x"C7",x"D1",x"D2",x"C7",x"CE",x"CE",x"D0",x"C8",x"CE",x"C7",x"C8",x"D6",x"00",x"02",x"50",x"54",x"D0",x"CF",x"C5",x"CE",x"D2",x"C8",x"C5",x"CF",x"D1",x"D0",x"CB",x"CA",x"03",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"01",x"4D",x"52",x"50",x"49",x"55",x"47",x"54",x"4E",x"4D",x"50",x"CD",x"CB",x"CD",x"C9",x"CF",x"D2",x"C7",x"D1",x"D0",x"CD",x"CD",x"C9",x"CF",x"00",x"3F",x"CA",x"CC",x"D1",x"CF",x"CF",x"C6",x"01",x"4C",x"CD",x"CC",x"CD",x"CA",x"CD",x"CC",x"00",x"52",x"4D",x"4D",x"50",x"4F",x"51",x"4D",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E"),
		(x"00",x"CD",x"4C",x"4F",x"4F",x"4F",x"4E",x"4F",x"54",x"53",x"50",x"00",x"CF",x"D1",x"C7",x"D1",x"CD",x"CC",x"D2",x"C6",x"CD",x"CE",x"00",x"02",x"01",x"53",x"48",x"01",x"CC",x"CE",x"C8",x"CF",x"D6",x"C9",x"C5",x"CB",x"CB",x"CD",x"00",x"00",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"4A",x"4F",x"4C",x"4C",x"4A",x"57",x"45",x"4B",x"56",x"45",x"01",x"CA",x"CD",x"C8",x"CC",x"C4",x"D1",x"CA",x"C6",x"CF",x"CB",x"CB",x"CC",x"02",x"56",x"CD",x"C7",x"CA",x"C6",x"D2",x"CF",x"00",x"56",x"C5",x"C7",x"C8",x"CC",x"D0",x"CD",x"02",x"50",x"48",x"4E",x"53",x"51",x"50",x"4F",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E"),
		(x"00",x"CD",x"4C",x"4F",x"4F",x"4F",x"4E",x"4F",x"4C",x"51",x"4C",x"07",x"CC",x"BC",x"CF",x"CA",x"CB",x"C9",x"C6",x"CD",x"C9",x"D1",x"00",x"00",x"02",x"44",x"54",x"01",x"C8",x"D1",x"C8",x"CC",x"C8",x"D3",x"C7",x"CD",x"C8",x"C9",x"02",x"00",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"05",x"57",x"4C",x"49",x"51",x"4C",x"4C",x"53",x"4F",x"4C",x"4C",x"05",x"CE",x"CB",x"CE",x"CE",x"CD",x"CC",x"CA",x"CB",x"C9",x"CF",x"C7",x"CD",x"01",x"55",x"C6",x"CC",x"D5",x"C4",x"CD",x"CB",x"07",x"49",x"D2",x"CD",x"CD",x"CE",x"CD",x"C9",x"01",x"52",x"4D",x"4F",x"50",x"53",x"50",x"4D",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E"),
		(x"00",x"CD",x"4C",x"4F",x"4F",x"4F",x"4E",x"4F",x"51",x"56",x"4E",x"55",x"08",x"C9",x"C7",x"CB",x"CA",x"CD",x"D2",x"BF",x"C6",x"06",x"03",x"00",x"51",x"56",x"4E",x"55",x"08",x"C9",x"C7",x"CB",x"CA",x"CD",x"D2",x"BF",x"C6",x"06",x"03",x"00",x"52",x"51",x"C4",x"CD",x"D8",x"CF",x"C4",x"C9",x"01",x"52",x"4D",x"4F",x"50",x"53",x"50",x"4D",x"51",x"56",x"4E",x"55",x"08",x"C9",x"C7",x"CB",x"CB",x"CB",x"CB",x"CB",x"CB",x"CB",x"CB",x"CB",x"00",x"53",x"CB",x"CF",x"C4",x"CD",x"D4",x"C4",x"00",x"53",x"CB",x"CF",x"C4",x"CD",x"D4",x"C4",x"01",x"52",x"4D",x"4F",x"50",x"53",x"50",x"4D",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E"),
		(x"00",x"CD",x"4C",x"4F",x"4F",x"4F",x"4E",x"4F",x"4C",x"47",x"4B",x"47",x"00",x"05",x"08",x"04",x"01",x"04",x"00",x"00",x"00",x"03",x"02",x"00",x"4C",x"47",x"4B",x"47",x"00",x"05",x"08",x"04",x"01",x"04",x"00",x"00",x"00",x"03",x"02",x"00",x"46",x"53",x"52",x"00",x"00",x"01",x"00",x"03",x"02",x"50",x"48",x"4E",x"53",x"51",x"50",x"4F",x"4C",x"47",x"4B",x"47",x"00",x"05",x"08",x"04",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"4B",x"4F",x"00",x"00",x"08",x"06",x"00",x"00",x"4B",x"4F",x"00",x"00",x"08",x"06",x"00",x"02",x"50",x"48",x"4E",x"53",x"51",x"50",x"4F",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E"),
		(x"00",x"CD",x"4C",x"4F",x"4F",x"4F",x"4E",x"4F",x"50",x"4C",x"50",x"55",x"4A",x"00",x"00",x"10",x"00",x"0B",x"03",x"06",x"02",x"00",x"00",x"4F",x"50",x"4C",x"50",x"55",x"4A",x"00",x"00",x"10",x"00",x"0B",x"03",x"06",x"02",x"00",x"00",x"4F",x"4B",x"53",x"4C",x"00",x"01",x"00",x"00",x"05",x"00",x"52",x"4D",x"4D",x"50",x"4F",x"51",x"4D",x"50",x"4C",x"50",x"55",x"4A",x"00",x"00",x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"4B",x"57",x"07",x"02",x"00",x"06",x"02",x"08",x"4B",x"57",x"07",x"02",x"00",x"06",x"02",x"00",x"52",x"4D",x"4D",x"50",x"4F",x"51",x"4D",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E"),
		(x"00",x"CD",x"4C",x"4F",x"4F",x"4F",x"4E",x"4F",x"54",x"4E",x"4F",x"4E",x"4B",x"00",x"00",x"00",x"03",x"00",x"00",x"06",x"00",x"04",x"04",x"4D",x"54",x"4E",x"4F",x"4E",x"4B",x"00",x"00",x"00",x"03",x"00",x"00",x"06",x"00",x"04",x"04",x"4D",x"4C",x"4F",x"57",x"00",x"00",x"01",x"00",x"04",x"00",x"56",x"56",x"4C",x"4B",x"4D",x"52",x"4C",x"54",x"4E",x"4F",x"4E",x"4B",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"4B",x"4A",x"00",x"01",x"00",x"05",x"03",x"00",x"4B",x"4A",x"00",x"01",x"00",x"05",x"03",x"00",x"56",x"56",x"4C",x"4B",x"4D",x"52",x"4C",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E"),
		(x"00",x"CD",x"4C",x"4F",x"4F",x"4F",x"4E",x"4F",x"49",x"50",x"4F",x"55",x"4C",x"52",x"00",x"03",x"03",x"02",x"00",x"00",x"08",x"00",x"4D",x"54",x"49",x"50",x"4F",x"55",x"4C",x"52",x"00",x"03",x"03",x"02",x"00",x"00",x"08",x"00",x"4D",x"54",x"50",x"5A",x"4A",x"04",x"01",x"00",x"00",x"03",x"00",x"42",x"4C",x"4C",x"51",x"50",x"50",x"4A",x"49",x"50",x"4F",x"55",x"4C",x"52",x"00",x"03",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"59",x"55",x"00",x"00",x"05",x"04",x"00",x"00",x"59",x"55",x"00",x"00",x"05",x"04",x"00",x"00",x"42",x"4C",x"4C",x"51",x"50",x"50",x"4A",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E"),
		(x"00",x"CD",x"4C",x"4F",x"4F",x"4F",x"4E",x"4F",x"50",x"4C",x"50",x"50",x"4F",x"45",x"54",x"48",x"53",x"53",x"4C",x"4E",x"4D",x"54",x"43",x"4D",x"50",x"4C",x"50",x"50",x"4F",x"45",x"54",x"48",x"53",x"53",x"4C",x"4E",x"4D",x"54",x"43",x"4D",x"4B",x"4F",x"45",x"54",x"55",x"4D",x"4E",x"50",x"53",x"5E",x"53",x"4B",x"4B",x"4A",x"4C",x"54",x"50",x"4C",x"50",x"50",x"4F",x"45",x"54",x"48",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"59",x"49",x"4A",x"49",x"51",x"4B",x"50",x"4A",x"59",x"49",x"4A",x"49",x"51",x"4B",x"50",x"4A",x"53",x"5E",x"53",x"4B",x"4B",x"4A",x"4C",x"54",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E"),
		(x"00",x"CD",x"4C",x"4F",x"4F",x"4F",x"4E",x"4F",x"52",x"4F",x"4D",x"4E",x"52",x"4A",x"4F",x"57",x"4E",x"4C",x"53",x"53",x"4C",x"53",x"50",x"47",x"52",x"4F",x"4D",x"4E",x"52",x"4A",x"4F",x"57",x"4E",x"4C",x"53",x"53",x"4C",x"53",x"50",x"47",x"51",x"4C",x"49",x"57",x"4C",x"52",x"57",x"48",x"4D",x"47",x"50",x"50",x"52",x"53",x"48",x"4C",x"52",x"4F",x"4D",x"4E",x"52",x"4A",x"4F",x"57",x"4C",x"4C",x"4C",x"4C",x"4C",x"4C",x"4C",x"4C",x"4E",x"4C",x"54",x"4D",x"50",x"55",x"4F",x"47",x"4E",x"4C",x"54",x"4D",x"50",x"55",x"4F",x"47",x"4D",x"47",x"50",x"50",x"52",x"53",x"48",x"4C",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E"),
		(x"00",x"CD",x"4C",x"4F",x"4F",x"4F",x"4E",x"4F",x"4C",x"4B",x"4F",x"54",x"4C",x"4E",x"4E",x"50",x"4D",x"4E",x"4D",x"53",x"4C",x"48",x"4B",x"58",x"4C",x"4B",x"4F",x"54",x"4C",x"4E",x"4E",x"50",x"4D",x"4E",x"4D",x"53",x"4C",x"48",x"4B",x"58",x"4F",x"4D",x"57",x"43",x"4F",x"53",x"46",x"51",x"52",x"48",x"58",x"4A",x"47",x"54",x"4D",x"4F",x"4C",x"4B",x"4F",x"54",x"4C",x"4E",x"4E",x"50",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"51",x"50",x"49",x"54",x"52",x"4B",x"4C",x"4B",x"57",x"50",x"49",x"54",x"52",x"4B",x"4C",x"4B",x"57",x"52",x"48",x"58",x"4A",x"47",x"54",x"4D",x"4F",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E"),
		(x"00",x"CD",x"4C",x"4F",x"4F",x"4F",x"4E",x"4F",x"4F",x"47",x"51",x"4F",x"51",x"4C",x"52",x"53",x"55",x"4B",x"54",x"51",x"44",x"4B",x"4E",x"4C",x"4C",x"54",x"4D",x"4C",x"4F",x"50",x"4D",x"4D",x"4F",x"47",x"51",x"4F",x"51",x"4C",x"52",x"53",x"4C",x"54",x"4D",x"4C",x"4F",x"50",x"4D",x"4D",x"4B",x"4A",x"51",x"51",x"4C",x"4F",x"49",x"49",x"4C",x"54",x"4D",x"4C",x"4F",x"50",x"4D",x"4D",x"4B",x"4A",x"51",x"51",x"4C",x"4F",x"49",x"49",x"50",x"4D",x"4A",x"4C",x"50",x"52",x"54",x"47",x"4C",x"54",x"4D",x"4C",x"4F",x"50",x"4D",x"4D",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4B",x"4A",x"51",x"51",x"4C",x"4F",x"49",x"49",x"4C",x"54",x"4D",x"4C",x"4F",x"50",x"4D",x"4D",x"4B",x"4A",x"51",x"51",x"4C",x"4F",x"49",x"49",x"4C",x"54",x"4D",x"4C",x"4F",x"50",x"4D",x"4D",x"4F",x"47",x"51",x"4F",x"51",x"4C",x"52",x"53",x"4C",x"54",x"4D",x"4C",x"4F",x"50",x"4D",x"4D",x"4F",x"47",x"51",x"4F",x"51",x"4C",x"52",x"53",x"4C",x"54",x"4D",x"4C",x"4F",x"50",x"4D",x"4D",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E"),
		(x"00",x"CD",x"4C",x"4F",x"4F",x"4F",x"4E",x"4F",x"50",x"4C",x"4E",x"4B",x"55",x"C9",x"C9",x"C0",x"C6",x"CD",x"4A",x"52",x"54",x"51",x"56",x"53",x"D2",x"C6",x"C6",x"CA",x"C6",x"50",x"54",x"4A",x"50",x"4C",x"4E",x"4B",x"55",x"C9",x"C9",x"C0",x"D2",x"C6",x"C6",x"CA",x"C6",x"50",x"54",x"4A",x"4E",x"58",x"C7",x"C8",x"D1",x"D0",x"C7",x"D0",x"D2",x"C6",x"C6",x"CA",x"C6",x"50",x"54",x"4A",x"4E",x"58",x"C7",x"C8",x"D1",x"D0",x"C7",x"D0",x"4F",x"50",x"50",x"4D",x"54",x"C4",x"C8",x"D3",x"D2",x"C6",x"C6",x"CA",x"C6",x"50",x"54",x"4A",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"58",x"C7",x"C8",x"D1",x"D0",x"C7",x"D0",x"D2",x"C6",x"C6",x"CA",x"C6",x"50",x"54",x"4A",x"4E",x"58",x"C7",x"C8",x"D1",x"D0",x"C7",x"D0",x"D2",x"C6",x"C6",x"CA",x"C6",x"50",x"54",x"4A",x"50",x"4C",x"4E",x"4B",x"55",x"C9",x"C9",x"C0",x"D2",x"C6",x"C6",x"CA",x"C6",x"50",x"54",x"4A",x"50",x"4C",x"4E",x"4B",x"55",x"C9",x"C9",x"C0",x"D2",x"C6",x"C6",x"CA",x"C6",x"50",x"54",x"4A",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E"),
		(x"00",x"CD",x"4C",x"4F",x"4F",x"4F",x"4E",x"4F",x"4F",x"4F",x"40",x"53",x"C8",x"CE",x"C7",x"D2",x"C9",x"C7",x"CC",x"52",x"49",x"47",x"54",x"C7",x"C6",x"CE",x"D9",x"CA",x"CA",x"D0",x"50",x"54",x"4F",x"4F",x"40",x"53",x"C8",x"CE",x"C7",x"D2",x"C6",x"CE",x"D9",x"CA",x"CA",x"D0",x"50",x"54",x"53",x"4B",x"DB",x"CB",x"CD",x"CC",x"C9",x"D0",x"C6",x"CE",x"D9",x"CA",x"CA",x"D0",x"50",x"54",x"53",x"4B",x"DB",x"CB",x"CD",x"CC",x"C9",x"D0",x"58",x"51",x"4D",x"56",x"C2",x"D2",x"CB",x"D1",x"C6",x"CE",x"D9",x"CA",x"CA",x"D0",x"50",x"54",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"53",x"4B",x"DB",x"CB",x"CD",x"CC",x"C9",x"D0",x"C6",x"CE",x"D9",x"CA",x"CA",x"D0",x"50",x"54",x"53",x"4B",x"DB",x"CB",x"CD",x"CC",x"C9",x"D0",x"C6",x"CE",x"D9",x"CA",x"CA",x"D0",x"50",x"54",x"4F",x"4F",x"40",x"53",x"C8",x"CE",x"C7",x"D2",x"C6",x"CE",x"D9",x"CA",x"CA",x"D0",x"50",x"54",x"4F",x"4F",x"40",x"53",x"C8",x"CE",x"C7",x"D2",x"C6",x"CE",x"D9",x"CA",x"CA",x"D0",x"50",x"54",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E"),
		(x"00",x"CD",x"4C",x"4F",x"4F",x"4F",x"4E",x"4F",x"54",x"48",x"4F",x"4F",x"CB",x"D4",x"D9",x"C8",x"CC",x"CC",x"D2",x"4E",x"56",x"52",x"4C",x"CC",x"D3",x"CB",x"CA",x"D4",x"CA",x"C8",x"4F",x"49",x"54",x"48",x"4F",x"4F",x"CB",x"D4",x"D9",x"C8",x"D3",x"CB",x"CA",x"D4",x"CA",x"C8",x"4F",x"49",x"4A",x"48",x"C4",x"C7",x"C6",x"CC",x"D0",x"D1",x"D3",x"CB",x"CA",x"D4",x"CA",x"C8",x"4F",x"49",x"4A",x"48",x"C4",x"C7",x"C6",x"CC",x"D0",x"D1",x"4A",x"41",x"4D",x"50",x"D5",x"CA",x"C3",x"CF",x"D3",x"CB",x"CA",x"D4",x"CA",x"C8",x"4F",x"49",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4A",x"48",x"C4",x"C7",x"C6",x"CC",x"D0",x"D1",x"D3",x"CB",x"CA",x"D4",x"CA",x"C8",x"4F",x"49",x"4A",x"48",x"C4",x"C7",x"C6",x"CC",x"D0",x"D1",x"D3",x"CB",x"CA",x"D4",x"CA",x"C8",x"4F",x"49",x"54",x"48",x"4F",x"4F",x"CB",x"D4",x"D9",x"C8",x"D3",x"CB",x"CA",x"D4",x"CA",x"C8",x"4F",x"49",x"54",x"48",x"4F",x"4F",x"CB",x"D4",x"D9",x"C8",x"D3",x"CB",x"CA",x"D4",x"CA",x"C8",x"4F",x"49",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E"),
		(x"00",x"CD",x"4C",x"4F",x"4F",x"4F",x"4E",x"4F",x"52",x"47",x"57",x"C6",x"C9",x"D2",x"C9",x"CB",x"CA",x"D1",x"CC",x"C5",x"4F",x"4A",x"C4",x"CE",x"C7",x"CB",x"C4",x"C4",x"C9",x"C4",x"C6",x"50",x"52",x"47",x"57",x"C6",x"C9",x"D2",x"C9",x"CB",x"C7",x"CB",x"C4",x"C4",x"C9",x"C4",x"C6",x"50",x"47",x"56",x"C7",x"D1",x"CD",x"C9",x"C9",x"CB",x"C7",x"CB",x"C4",x"C4",x"C9",x"C4",x"C6",x"50",x"47",x"56",x"C7",x"D1",x"CD",x"C9",x"C9",x"CB",x"5C",x"4A",x"53",x"C5",x"CA",x"D1",x"C6",x"C9",x"C7",x"CB",x"C4",x"C4",x"C9",x"C4",x"C6",x"50",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"47",x"56",x"C7",x"D1",x"CD",x"C9",x"C9",x"CB",x"C7",x"CB",x"C4",x"C4",x"C9",x"C4",x"C6",x"50",x"47",x"56",x"C7",x"D1",x"CD",x"C9",x"C9",x"CB",x"C7",x"CB",x"C4",x"C4",x"C9",x"C4",x"C6",x"50",x"52",x"47",x"57",x"C6",x"C9",x"D2",x"C9",x"CB",x"C7",x"CB",x"C4",x"C4",x"C9",x"C4",x"C6",x"50",x"52",x"47",x"57",x"C6",x"C9",x"D2",x"C9",x"CB",x"C7",x"CB",x"C4",x"C4",x"C9",x"C4",x"C6",x"50",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E"),
		(x"00",x"CD",x"4C",x"4F",x"4F",x"4F",x"4E",x"4F",x"4F",x"4F",x"53",x"C4",x"C9",x"CB",x"CA",x"C6",x"CE",x"CA",x"CD",x"CB",x"50",x"52",x"CD",x"CC",x"CC",x"C6",x"D0",x"D1",x"CF",x"D4",x"C8",x"5B",x"4F",x"4F",x"53",x"C4",x"C9",x"CB",x"CA",x"C6",x"CC",x"C6",x"D0",x"D1",x"CF",x"D4",x"C8",x"5B",x"52",x"57",x"D1",x"CA",x"D1",x"CE",x"C8",x"D2",x"CC",x"C6",x"D0",x"D1",x"CF",x"D4",x"C8",x"5B",x"52",x"57",x"D1",x"CA",x"D1",x"CE",x"C8",x"D2",x"00",x"4D",x"63",x"CA",x"C8",x"CA",x"CA",x"CB",x"CC",x"C6",x"D0",x"D1",x"CF",x"D4",x"C8",x"5B",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"52",x"57",x"D1",x"CA",x"D1",x"CE",x"C8",x"D2",x"CC",x"C6",x"D0",x"D1",x"CF",x"D4",x"C8",x"5B",x"52",x"57",x"D1",x"CA",x"D1",x"CE",x"C8",x"D2",x"CC",x"C6",x"D0",x"D1",x"CF",x"D4",x"C8",x"5B",x"4F",x"4F",x"53",x"C4",x"C9",x"CB",x"CA",x"C6",x"CC",x"C6",x"D0",x"D1",x"CF",x"D4",x"C8",x"5B",x"4F",x"4F",x"53",x"C4",x"C9",x"CB",x"CA",x"C6",x"CC",x"C6",x"D0",x"D1",x"CF",x"D4",x"C8",x"5B",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E"),
		(x"00",x"CD",x"4C",x"4F",x"4F",x"4F",x"4E",x"4F",x"4E",x"54",x"CB",x"CA",x"CF",x"C9",x"D0",x"CD",x"CB",x"CF",x"C9",x"D1",x"C3",x"CB",x"C8",x"CD",x"CD",x"CC",x"CD",x"CC",x"CE",x"C7",x"CF",x"CB",x"4E",x"54",x"CB",x"CA",x"CF",x"C9",x"D0",x"CD",x"CD",x"CC",x"CD",x"CC",x"CE",x"C7",x"CF",x"CB",x"4F",x"4C",x"CD",x"C6",x"CE",x"CD",x"C5",x"C9",x"CD",x"CC",x"CD",x"CC",x"CE",x"C7",x"CF",x"CB",x"4F",x"4C",x"CD",x"C6",x"CE",x"CD",x"C5",x"C9",x"07",x"49",x"C5",x"D1",x"C6",x"CB",x"DA",x"CD",x"CD",x"CC",x"CD",x"CC",x"CE",x"C7",x"CF",x"CB",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4F",x"4C",x"CD",x"C6",x"CE",x"CD",x"C5",x"C9",x"CD",x"CC",x"CD",x"CC",x"CE",x"C7",x"CF",x"CB",x"4F",x"4C",x"CD",x"C6",x"CE",x"CD",x"C5",x"C9",x"CD",x"CC",x"CD",x"CC",x"CE",x"C7",x"CF",x"CB",x"4E",x"54",x"CB",x"CA",x"CF",x"C9",x"D0",x"CD",x"CD",x"CC",x"CD",x"CC",x"CE",x"C7",x"CF",x"CB",x"4E",x"54",x"CB",x"CA",x"CF",x"C9",x"D0",x"CD",x"CD",x"CC",x"CD",x"CC",x"CE",x"C7",x"CF",x"CB",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E"),
		(x"00",x"CD",x"4C",x"4F",x"4F",x"4F",x"4E",x"4F",x"47",x"52",x"CE",x"C7",x"CE",x"C8",x"C6",x"D2",x"CE",x"CB",x"CD",x"C0",x"D7",x"D1",x"C7",x"CC",x"CC",x"D2",x"C6",x"CB",x"CB",x"CE",x"C8",x"CB",x"47",x"52",x"CE",x"C7",x"CE",x"C8",x"C6",x"D2",x"CC",x"D2",x"C6",x"CB",x"CB",x"CE",x"C8",x"CB",x"4C",x"52",x"CA",x"CF",x"C9",x"CA",x"CE",x"CF",x"CC",x"D2",x"C6",x"CB",x"CB",x"CE",x"C8",x"CB",x"4C",x"52",x"CA",x"CF",x"C9",x"CA",x"CE",x"CF",x"02",x"50",x"CA",x"CE",x"C7",x"CF",x"CA",x"C5",x"CC",x"D2",x"C6",x"CB",x"CB",x"CE",x"C8",x"CB",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4C",x"52",x"CA",x"CF",x"C9",x"CA",x"CE",x"CF",x"CC",x"D2",x"C6",x"CB",x"CB",x"CE",x"C8",x"CB",x"4C",x"52",x"CA",x"CF",x"C9",x"CA",x"CE",x"CF",x"CC",x"D2",x"C6",x"CB",x"CB",x"CE",x"C8",x"CB",x"47",x"52",x"CE",x"C7",x"CE",x"C8",x"C6",x"D2",x"CC",x"D2",x"C6",x"CB",x"CB",x"CE",x"C8",x"CB",x"47",x"52",x"CE",x"C7",x"CE",x"C8",x"C6",x"D2",x"CC",x"D2",x"C6",x"CB",x"CB",x"CE",x"C8",x"CB",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E"),
		(x"00",x"CD",x"4C",x"4F",x"4F",x"4F",x"4E",x"4F",x"4E",x"4E",x"CB",x"CE",x"C8",x"CD",x"CA",x"CC",x"D0",x"D5",x"C7",x"C9",x"CB",x"D2",x"C8",x"CF",x"D0",x"D5",x"C7",x"C9",x"CB",x"D2",x"C8",x"CF",x"53",x"50",x"C6",x"CF",x"CC",x"CD",x"CA",x"CE",x"D0",x"D5",x"C7",x"C9",x"CB",x"D2",x"C8",x"CF",x"53",x"50",x"C6",x"CF",x"CC",x"CD",x"CA",x"CE",x"D0",x"D5",x"C7",x"C9",x"CB",x"D2",x"C8",x"CF",x"53",x"50",x"C6",x"CF",x"CC",x"CD",x"CA",x"CE",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"D0",x"D5",x"C7",x"C9",x"CB",x"D2",x"C8",x"CF",x"53",x"4E",x"4A",x"52",x"4D",x"51",x"4D",x"51",x"4E",x"4E",x"CB",x"CE",x"C8",x"CD",x"CA",x"CC",x"D0",x"D5",x"C7",x"C9",x"CB",x"D2",x"C8",x"CF",x"53",x"50",x"C6",x"CF",x"CC",x"CD",x"CA",x"CE",x"D0",x"D5",x"C7",x"C9",x"CB",x"D2",x"C8",x"CF",x"53",x"50",x"C6",x"CF",x"CC",x"CD",x"CA",x"CE",x"D0",x"D5",x"C7",x"C9",x"CB",x"D2",x"C8",x"CF",x"53",x"50",x"C6",x"CF",x"CC",x"CD",x"CA",x"CE",x"D0",x"D5",x"C7",x"C9",x"CB",x"D2",x"C8",x"CF",x"53",x"4E",x"4A",x"52",x"4D",x"51",x"4D",x"51",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E"),
		(x"00",x"CD",x"4C",x"4F",x"4F",x"4F",x"4E",x"4F",x"4E",x"4E",x"CB",x"CE",x"C8",x"CD",x"CA",x"CC",x"00",x"00",x"CF",x"CB",x"CA",x"CB",x"CB",x"C4",x"00",x"00",x"CF",x"CB",x"CA",x"CB",x"CB",x"C4",x"00",x"41",x"CF",x"CD",x"C9",x"CF",x"CC",x"C8",x"00",x"00",x"CF",x"CB",x"CA",x"CB",x"CB",x"C4",x"00",x"41",x"CF",x"CD",x"C9",x"CF",x"CC",x"C8",x"00",x"00",x"CF",x"CB",x"CA",x"CB",x"CB",x"C4",x"00",x"41",x"CF",x"CD",x"C9",x"CF",x"CC",x"C8",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"00",x"CF",x"CB",x"CA",x"CB",x"CB",x"C4",x"00",x"40",x"52",x"50",x"4B",x"53",x"4E",x"4C",x"4E",x"4E",x"CB",x"CE",x"C8",x"CD",x"CA",x"CC",x"00",x"00",x"CF",x"CB",x"CA",x"CB",x"CB",x"C4",x"00",x"41",x"CF",x"CD",x"C9",x"CF",x"CC",x"C8",x"00",x"00",x"CF",x"CB",x"CA",x"CB",x"CB",x"C4",x"00",x"41",x"CF",x"CD",x"C9",x"CF",x"CC",x"C8",x"00",x"00",x"CF",x"CB",x"CA",x"CB",x"CB",x"C4",x"00",x"41",x"CF",x"CD",x"C9",x"CF",x"CC",x"C8",x"00",x"00",x"CF",x"CB",x"CA",x"CB",x"CB",x"C4",x"00",x"40",x"52",x"50",x"4B",x"53",x"4E",x"4C",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E"),
		(x"00",x"CD",x"4C",x"4F",x"4F",x"4F",x"4E",x"4F",x"4E",x"4E",x"CB",x"CE",x"C8",x"CD",x"CA",x"CC",x"00",x"0A",x"CA",x"D0",x"CD",x"C6",x"CC",x"D1",x"00",x"0A",x"CA",x"D0",x"CD",x"C6",x"CC",x"D1",x"00",x"51",x"D2",x"C9",x"C9",x"C8",x"C8",x"CE",x"00",x"0A",x"CA",x"D0",x"CD",x"C6",x"CC",x"D1",x"00",x"51",x"D2",x"C9",x"C9",x"C8",x"C8",x"CE",x"00",x"0A",x"CA",x"D0",x"CD",x"C6",x"CC",x"D1",x"00",x"51",x"D2",x"C9",x"C9",x"C8",x"C8",x"CE",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"0A",x"CA",x"D0",x"CD",x"C6",x"CC",x"D1",x"00",x"4F",x"56",x"4C",x"4B",x"4D",x"4B",x"52",x"4E",x"4E",x"CB",x"CE",x"C8",x"CD",x"CA",x"CC",x"00",x"0A",x"CA",x"D0",x"CD",x"C6",x"CC",x"D1",x"00",x"51",x"D2",x"C9",x"C9",x"C8",x"C8",x"CE",x"00",x"0A",x"CA",x"D0",x"CD",x"C6",x"CC",x"D1",x"00",x"51",x"D2",x"C9",x"C9",x"C8",x"C8",x"CE",x"00",x"0A",x"CA",x"D0",x"CD",x"C6",x"CC",x"D1",x"00",x"51",x"D2",x"C9",x"C9",x"C8",x"C8",x"CE",x"00",x"0A",x"CA",x"D0",x"CD",x"C6",x"CC",x"D1",x"00",x"4F",x"56",x"4C",x"4B",x"4D",x"4B",x"52",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E"),
		(x"00",x"CD",x"4C",x"4F",x"4F",x"4F",x"4E",x"4F",x"4E",x"4E",x"CB",x"CE",x"C8",x"CD",x"CA",x"CC",x"01",x"03",x"CB",x"CD",x"D3",x"C6",x"CA",x"CA",x"01",x"03",x"CB",x"CD",x"D3",x"C6",x"CA",x"CA",x"03",x"52",x"C8",x"CD",x"D2",x"C5",x"C7",x"CD",x"01",x"03",x"CB",x"CD",x"D3",x"C6",x"CA",x"CA",x"03",x"52",x"C8",x"CD",x"D2",x"C5",x"C7",x"CD",x"01",x"03",x"CB",x"CD",x"D3",x"C6",x"CA",x"CA",x"03",x"52",x"C8",x"CD",x"D2",x"C5",x"C7",x"CD",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"01",x"03",x"CB",x"CD",x"D3",x"C6",x"CA",x"CA",x"03",x"50",x"4D",x"4F",x"54",x"49",x"4A",x"50",x"4E",x"4E",x"CB",x"CE",x"C8",x"CD",x"CA",x"CC",x"01",x"03",x"CB",x"CD",x"D3",x"C6",x"CA",x"CA",x"03",x"52",x"C8",x"CD",x"D2",x"C5",x"C7",x"CD",x"01",x"03",x"CB",x"CD",x"D3",x"C6",x"CA",x"CA",x"03",x"52",x"C8",x"CD",x"D2",x"C5",x"C7",x"CD",x"01",x"03",x"CB",x"CD",x"D3",x"C6",x"CA",x"CA",x"03",x"52",x"C8",x"CD",x"D2",x"C5",x"C7",x"CD",x"01",x"03",x"CB",x"CD",x"D3",x"C6",x"CA",x"CA",x"03",x"50",x"4D",x"4F",x"54",x"49",x"4A",x"50",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E"),
		(x"00",x"CD",x"4C",x"4F",x"4F",x"4F",x"4E",x"4F",x"4E",x"4E",x"CB",x"CE",x"C8",x"CD",x"CA",x"CC",x"02",x"06",x"D0",x"C5",x"CF",x"C7",x"CC",x"CA",x"02",x"06",x"D0",x"C5",x"CF",x"C7",x"CC",x"CA",x"00",x"4D",x"CB",x"CC",x"CB",x"C8",x"D0",x"C8",x"02",x"06",x"D0",x"C5",x"CF",x"C7",x"CC",x"CA",x"00",x"4D",x"CB",x"CC",x"CB",x"C8",x"D0",x"C8",x"02",x"06",x"D0",x"C5",x"CF",x"C7",x"CC",x"CA",x"00",x"4D",x"CB",x"CC",x"CB",x"C8",x"D0",x"C8",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"02",x"06",x"D0",x"C5",x"CF",x"C7",x"CC",x"CA",x"00",x"4C",x"4E",x"4F",x"4D",x"4C",x"53",x"4C",x"4E",x"4E",x"CB",x"CE",x"C8",x"CD",x"CA",x"CC",x"02",x"06",x"D0",x"C5",x"CF",x"C7",x"CC",x"CA",x"00",x"4D",x"CB",x"CC",x"CB",x"C8",x"D0",x"C8",x"02",x"06",x"D0",x"C5",x"CF",x"C7",x"CC",x"CA",x"00",x"4D",x"CB",x"CC",x"CB",x"C8",x"D0",x"C8",x"02",x"06",x"D0",x"C5",x"CF",x"C7",x"CC",x"CA",x"00",x"4D",x"CB",x"CC",x"CB",x"C8",x"D0",x"C8",x"02",x"06",x"D0",x"C5",x"CF",x"C7",x"CC",x"CA",x"00",x"4C",x"4E",x"4F",x"4D",x"4C",x"53",x"4C",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E"),
		(x"00",x"CD",x"4C",x"4F",x"4F",x"4F",x"4E",x"4F",x"4E",x"4E",x"CB",x"CE",x"C8",x"CD",x"CA",x"CC",x"00",x"56",x"C0",x"C8",x"D2",x"CD",x"CB",x"CD",x"00",x"56",x"C0",x"C8",x"D2",x"CD",x"CB",x"CD",x"04",x"51",x"CD",x"CA",x"C6",x"C8",x"D4",x"C9",x"00",x"56",x"C0",x"C8",x"D2",x"CD",x"CB",x"CD",x"04",x"51",x"CD",x"CA",x"C6",x"C8",x"D4",x"C9",x"00",x"56",x"C0",x"C8",x"D2",x"CD",x"CB",x"CD",x"04",x"51",x"CD",x"CA",x"C6",x"C8",x"D4",x"C9",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"56",x"C0",x"C8",x"D2",x"CD",x"CB",x"CD",x"04",x"4F",x"51",x"4E",x"49",x"4C",x"56",x"4C",x"4E",x"4E",x"CB",x"CE",x"C8",x"CD",x"CA",x"CC",x"00",x"56",x"C0",x"C8",x"D2",x"CD",x"CB",x"CD",x"04",x"51",x"CD",x"CA",x"C6",x"C8",x"D4",x"C9",x"00",x"56",x"C0",x"C8",x"D2",x"CD",x"CB",x"CD",x"04",x"51",x"CD",x"CA",x"C6",x"C8",x"D4",x"C9",x"00",x"56",x"C0",x"C8",x"D2",x"CD",x"CB",x"CD",x"04",x"51",x"CD",x"CA",x"C6",x"C8",x"D4",x"C9",x"00",x"56",x"C0",x"C8",x"D2",x"CD",x"CB",x"CD",x"04",x"4F",x"51",x"4E",x"49",x"4C",x"56",x"4C",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E"),
		(x"00",x"CD",x"4C",x"4F",x"4F",x"4F",x"4E",x"4F",x"4E",x"4E",x"CB",x"CE",x"C8",x"CD",x"CA",x"CC",x"01",x"56",x"CE",x"C6",x"C7",x"C6",x"CB",x"CF",x"01",x"56",x"CE",x"C6",x"C7",x"C6",x"CB",x"CF",x"01",x"47",x"C7",x"CD",x"D1",x"CC",x"CC",x"C8",x"01",x"56",x"CE",x"C6",x"C7",x"C6",x"CB",x"CF",x"01",x"47",x"C7",x"CD",x"D1",x"CC",x"CC",x"C8",x"01",x"56",x"CE",x"C6",x"C7",x"C6",x"CB",x"CF",x"01",x"47",x"C7",x"CD",x"D1",x"CC",x"CC",x"C8",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"01",x"56",x"CE",x"C6",x"C7",x"C6",x"CB",x"CF",x"01",x"46",x"4B",x"50",x"53",x"4F",x"4E",x"4C",x"4E",x"4E",x"CB",x"CE",x"C8",x"CD",x"CA",x"CC",x"01",x"56",x"CE",x"C6",x"C7",x"C6",x"CB",x"CF",x"01",x"47",x"C7",x"CD",x"D1",x"CC",x"CC",x"C8",x"01",x"56",x"CE",x"C6",x"C7",x"C6",x"CB",x"CF",x"01",x"47",x"C7",x"CD",x"D1",x"CC",x"CC",x"C8",x"01",x"56",x"CE",x"C6",x"C7",x"C6",x"CB",x"CF",x"01",x"47",x"C7",x"CD",x"D1",x"CC",x"CC",x"C8",x"01",x"56",x"CE",x"C6",x"C7",x"C6",x"CB",x"CF",x"01",x"46",x"4B",x"50",x"53",x"4F",x"4E",x"4C",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E"),
		(x"00",x"CD",x"4C",x"4F",x"4F",x"4F",x"4E",x"4F",x"4E",x"4E",x"CB",x"CE",x"C8",x"CD",x"CA",x"CC",x"03",x"47",x"CB",x"C8",x"D1",x"CF",x"CA",x"CC",x"03",x"47",x"CB",x"C8",x"D1",x"CF",x"CA",x"CC",x"02",x"51",x"CF",x"C9",x"CE",x"CA",x"C8",x"CD",x"03",x"47",x"CB",x"C8",x"D1",x"CF",x"CA",x"CC",x"02",x"51",x"CF",x"C9",x"CE",x"CA",x"C8",x"CD",x"03",x"47",x"CB",x"C8",x"D1",x"CF",x"CA",x"CC",x"02",x"51",x"CF",x"C9",x"CE",x"CA",x"C8",x"CD",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"03",x"47",x"CB",x"C8",x"D1",x"CF",x"CA",x"CC",x"02",x"50",x"53",x"4D",x"4F",x"4E",x"4A",x"51",x"4E",x"4E",x"CB",x"CE",x"C8",x"CD",x"CA",x"CC",x"03",x"47",x"CB",x"C8",x"D1",x"CF",x"CA",x"CC",x"02",x"51",x"CF",x"C9",x"CE",x"CA",x"C8",x"CD",x"03",x"47",x"CB",x"C8",x"D1",x"CF",x"CA",x"CC",x"02",x"51",x"CF",x"C9",x"CE",x"CA",x"C8",x"CD",x"03",x"47",x"CB",x"C8",x"D1",x"CF",x"CA",x"CC",x"02",x"51",x"CF",x"C9",x"CE",x"CA",x"C8",x"CD",x"03",x"47",x"CB",x"C8",x"D1",x"CF",x"CA",x"CC",x"02",x"50",x"53",x"4D",x"4F",x"4E",x"4A",x"51",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E"),
		(x"00",x"CD",x"4C",x"4F",x"4F",x"4F",x"4E",x"4F",x"4E",x"4E",x"CB",x"CE",x"C8",x"CD",x"CA",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"04",x"4D",x"CA",x"C8",x"CD",x"CA",x"CF",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"4D",x"50",x"4E",x"4E",x"4E",x"50",x"4D",x"4E",x"4E",x"CB",x"CE",x"C8",x"CD",x"CA",x"CC",x"04",x"4D",x"CA",x"C8",x"CD",x"CA",x"CF",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"04",x"4D",x"CA",x"C8",x"CD",x"CA",x"CF",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"52",x"CB",x"CD",x"CA",x"C7",x"CE",x"CD",x"01",x"4A",x"D1",x"CC",x"CD",x"D0",x"CA",x"D4",x"01",x"52",x"4D",x"4F",x"50",x"53",x"50",x"4D",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E"),
		(x"00",x"CD",x"4C",x"4F",x"4F",x"4F",x"4E",x"4F",x"4E",x"4E",x"CB",x"CE",x"C8",x"CD",x"CA",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"CF",x"C8",x"D0",x"D0",x"CF",x"C8",x"CA",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"4D",x"50",x"4E",x"4E",x"4E",x"50",x"4D",x"4E",x"4E",x"CB",x"CE",x"C8",x"CD",x"CA",x"CC",x"00",x"CF",x"C8",x"D0",x"D0",x"CF",x"C8",x"CA",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"CF",x"C8",x"D0",x"D0",x"CF",x"C8",x"CA",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"05",x"57",x"C2",x"CE",x"CF",x"CC",x"C9",x"CA",x"C7",x"55",x"4B",x"00",x"00",x"01",x"04",x"00",x"02",x"50",x"48",x"4E",x"53",x"51",x"50",x"4F",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E"),
		(x"00",x"CD",x"4C",x"4F",x"4F",x"4F",x"4E",x"4F",x"4E",x"4E",x"CB",x"CE",x"C8",x"CD",x"CA",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"03",x"C5",x"CC",x"CA",x"D3",x"CD",x"C1",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"4D",x"50",x"4E",x"4E",x"4E",x"50",x"4D",x"4E",x"4E",x"CB",x"CE",x"C8",x"CD",x"CA",x"CC",x"03",x"C5",x"CC",x"CA",x"D3",x"CD",x"C1",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"03",x"C5",x"CC",x"CA",x"D3",x"CD",x"C1",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"01",x"56",x"C9",x"C5",x"D1",x"CD",x"CC",x"C8",x"CE",x"CE",x"58",x"05",x"00",x"06",x"01",x"03",x"00",x"52",x"4D",x"4D",x"50",x"4F",x"51",x"4D",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E"),
		(x"00",x"CD",x"4C",x"4F",x"4F",x"4F",x"4E",x"4F",x"4E",x"4E",x"CB",x"CE",x"C8",x"CD",x"CA",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"D4",x"C9",x"CC",x"CF",x"CC",x"D0",x"D1",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"4D",x"50",x"4E",x"4E",x"4E",x"50",x"4D",x"4E",x"4E",x"CB",x"CE",x"C8",x"CD",x"CA",x"CC",x"00",x"D4",x"C9",x"CC",x"CF",x"CC",x"D0",x"D1",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"D4",x"C9",x"CC",x"CF",x"CC",x"D0",x"D1",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"4A",x"51",x"CB",x"C7",x"CD",x"C9",x"D1",x"CC",x"C7",x"C9",x"D0",x"02",x"00",x"00",x"02",x"00",x"56",x"56",x"4C",x"4B",x"4D",x"52",x"4C",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E"),
		(x"00",x"CD",x"4C",x"4F",x"4F",x"4F",x"4E",x"4F",x"4E",x"4E",x"CB",x"CE",x"C8",x"CD",x"CA",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"08",x"C5",x"CA",x"D5",x"C5",x"CA",x"D1",x"01",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"4D",x"50",x"4E",x"4E",x"4E",x"50",x"4D",x"4E",x"4E",x"CB",x"CE",x"C8",x"CD",x"CA",x"CC",x"08",x"C5",x"CA",x"D5",x"C5",x"CA",x"D1",x"01",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"08",x"C5",x"CA",x"D5",x"C5",x"CA",x"D1",x"01",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"51",x"4C",x"C3",x"CF",x"CE",x"D2",x"CE",x"CB",x"C8",x"CD",x"C5",x"D2",x"CF",x"00",x"00",x"00",x"42",x"4C",x"4C",x"51",x"50",x"50",x"4A",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E"),
		(x"00",x"CD",x"4C",x"4F",x"4F",x"4F",x"4E",x"4F",x"4E",x"4E",x"CB",x"CE",x"C8",x"CD",x"CA",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"04",x"D0",x"C2",x"CD",x"C7",x"CE",x"00",x"01",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"4D",x"50",x"4E",x"4E",x"4E",x"50",x"4D",x"4E",x"4E",x"CB",x"CE",x"C8",x"CD",x"CA",x"CC",x"04",x"D0",x"C2",x"CD",x"C7",x"CE",x"00",x"01",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"04",x"D0",x"C2",x"CD",x"C7",x"CE",x"00",x"01",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"03",x"4D",x"55",x"00",x"C9",x"D8",x"C2",x"BE",x"D0",x"C6",x"C3",x"D9",x"CE",x"C8",x"CE",x"53",x"53",x"5E",x"53",x"4B",x"4B",x"4A",x"4C",x"54",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E"),
		(x"00",x"CD",x"4C",x"4F",x"4F",x"4F",x"4E",x"4F",x"4E",x"4E",x"CB",x"CE",x"C8",x"CD",x"CA",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"D0",x"C9",x"D2",x"C8",x"C6",x"D1",x"00",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"4D",x"50",x"4E",x"4E",x"4E",x"50",x"4D",x"4E",x"4E",x"CB",x"CE",x"C8",x"CD",x"CA",x"CC",x"00",x"D0",x"C9",x"D2",x"C8",x"C6",x"D1",x"00",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"D0",x"C9",x"D2",x"C8",x"C6",x"D1",x"00",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"04",x"49",x"4F",x"00",x"00",x"00",x"D6",x"CC",x"CB",x"D2",x"C9",x"D1",x"C8",x"C5",x"CC",x"50",x"4D",x"47",x"50",x"50",x"52",x"53",x"48",x"4C",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E"),
		(x"00",x"CD",x"4C",x"4F",x"4F",x"4F",x"4E",x"4F",x"4E",x"4E",x"CB",x"CE",x"C8",x"CD",x"CA",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"01",x"C8",x"CD",x"D0",x"CD",x"CB",x"CB",x"CF",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"4D",x"50",x"4E",x"4E",x"4E",x"50",x"4D",x"4E",x"4E",x"CB",x"CE",x"C8",x"CD",x"CA",x"CC",x"01",x"C8",x"CD",x"D0",x"CD",x"CB",x"CB",x"CF",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"01",x"C8",x"CD",x"D0",x"CD",x"CB",x"CB",x"CF",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"05",x"47",x"52",x"4D",x"07",x"00",x"01",x"06",x"CB",x"CB",x"D0",x"C8",x"C6",x"D1",x"CC",x"CB",x"52",x"48",x"58",x"4A",x"47",x"54",x"4D",x"4F",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E"),
		(x"00",x"CD",x"4C",x"4F",x"4F",x"4F",x"4E",x"4F",x"4E",x"4E",x"CB",x"CE",x"C8",x"CD",x"CA",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"57",x"C9",x"C9",x"CB",x"C9",x"C8",x"CF",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"CF",x"C8",x"C9",x"CE",x"CF",x"C8",x"CE",x"54",x"46",x"D4",x"C8",x"C3",x"D0",x"CE",x"CB",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"4D",x"50",x"4E",x"4E",x"4E",x"50",x"4D",x"4E",x"4E",x"CB",x"CE",x"C8",x"CD",x"CA",x"CC",x"00",x"D0",x"C9",x"D0",x"C6",x"CF",x"CC",x"CC",x"54",x"46",x"D4",x"C8",x"C3",x"D0",x"CE",x"CB",x"00",x"CF",x"C8",x"C9",x"CE",x"CF",x"C8",x"CE",x"54",x"46",x"D4",x"C8",x"C3",x"D0",x"CE",x"CB",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"47",x"4D",x"54",x"00",x"03",x"03",x"00",x"00",x"02",x"CE",x"CE",x"C9",x"CD",x"D5",x"C2",x"52",x"48",x"58",x"4A",x"47",x"54",x"4D",x"4F",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E"),
		(x"00",x"CD",x"4C",x"4F",x"4F",x"4F",x"4E",x"4F",x"4E",x"4E",x"CB",x"CE",x"C8",x"CD",x"CA",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"CF",x"C8",x"D1",x"C4",x"D1",x"CE",x"C8",x"CE",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"55",x"CF",x"CA",x"CB",x"CE",x"C9",x"D0",x"4E",x"44",x"CC",x"CF",x"CE",x"CF",x"C9",x"C8",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"4D",x"50",x"4E",x"4E",x"4E",x"50",x"4D",x"4E",x"4E",x"CB",x"CE",x"C8",x"CD",x"CA",x"CC",x"00",x"00",x"C6",x"D3",x"CA",x"C7",x"CF",x"CB",x"4E",x"44",x"CC",x"CF",x"CE",x"CF",x"C9",x"C8",x"00",x"55",x"CF",x"CA",x"CB",x"CE",x"C9",x"D0",x"4E",x"44",x"CC",x"CF",x"CE",x"CF",x"C9",x"C8",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"0A",x"56",x"CA",x"CF",x"CE",x"D2",x"D1",x"C8",x"09",x"00",x"CA",x"CE",x"CC",x"D0",x"C8",x"D2",x"4D",x"47",x"50",x"50",x"52",x"53",x"48",x"4C",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E"),
		(x"00",x"CD",x"4C",x"4F",x"4F",x"4F",x"4E",x"4F",x"4E",x"4E",x"CB",x"CE",x"C8",x"CD",x"CA",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"D1",x"CC",x"CC",x"CB",x"CE",x"CB",x"C9",x"CD",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"07",x"41",x"D1",x"D2",x"C8",x"D0",x"C7",x"CB",x"54",x"5C",x"D1",x"CA",x"C7",x"C6",x"CB",x"D1",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"4D",x"50",x"4E",x"4E",x"4E",x"50",x"4D",x"4E",x"4E",x"CB",x"CE",x"C8",x"CD",x"CA",x"CC",x"04",x"03",x"CA",x"CD",x"C5",x"CE",x"CA",x"CA",x"54",x"5C",x"D1",x"CA",x"C7",x"C6",x"CB",x"D1",x"07",x"41",x"D1",x"D2",x"C8",x"D0",x"C7",x"CB",x"54",x"5C",x"D1",x"CA",x"C7",x"C6",x"CB",x"D1",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"47",x"D1",x"C3",x"CE",x"CD",x"C8",x"CE",x"00",x"00",x"C6",x"C4",x"CF",x"C8",x"D1",x"CF",x"53",x"5E",x"53",x"4B",x"4B",x"4A",x"4C",x"54",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E"),
		(x"00",x"CD",x"4C",x"4F",x"4F",x"4F",x"4E",x"4F",x"4E",x"4E",x"CB",x"CE",x"C8",x"CD",x"CA",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"C9",x"D2",x"CF",x"CD",x"C2",x"C9",x"CE",x"CE",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"58",x"C6",x"CF",x"C6",x"D1",x"C8",x"CC",x"00",x"40",x"CA",x"CB",x"CC",x"CC",x"CF",x"C6",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"4D",x"50",x"4E",x"4E",x"4E",x"50",x"4D",x"4E",x"4E",x"CB",x"CE",x"C8",x"CD",x"CA",x"CC",x"01",x"03",x"CF",x"CA",x"CB",x"CE",x"C8",x"CA",x"00",x"40",x"CA",x"CB",x"CC",x"CC",x"CF",x"C6",x"00",x"58",x"C6",x"CF",x"C6",x"D1",x"C8",x"CC",x"00",x"40",x"CA",x"CB",x"CC",x"CC",x"CF",x"C6",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"55",x"CA",x"CB",x"C8",x"C8",x"CB",x"D5",x"5B",x"01",x"D6",x"CD",x"D4",x"C8",x"C8",x"C7",x"00",x"42",x"4C",x"4C",x"51",x"50",x"50",x"4A",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E"),
		(x"00",x"CD",x"4C",x"4F",x"4F",x"4F",x"4E",x"4F",x"4E",x"4E",x"CB",x"CE",x"C8",x"CD",x"CA",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"CB",x"C8",x"C4",x"D3",x"CC",x"CF",x"CD",x"C9",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"48",x"CA",x"CD",x"CB",x"CC",x"CB",x"CD",x"00",x"53",x"D3",x"CB",x"C8",x"C9",x"D3",x"C8",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"4D",x"50",x"4E",x"4E",x"4E",x"50",x"4D",x"4E",x"4E",x"CB",x"CE",x"C8",x"CD",x"CA",x"CC",x"02",x"00",x"C9",x"CC",x"CD",x"C9",x"CF",x"C9",x"00",x"53",x"D3",x"CB",x"C8",x"C9",x"D3",x"C8",x"00",x"48",x"CA",x"CD",x"CB",x"CC",x"CB",x"CD",x"00",x"53",x"D3",x"CB",x"C8",x"C9",x"D3",x"C8",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"01",x"56",x"CA",x"CD",x"D0",x"C7",x"CD",x"C7",x"51",x"00",x"CF",x"CB",x"C5",x"C7",x"D7",x"C6",x"00",x"56",x"56",x"4C",x"4B",x"4D",x"52",x"4C",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E"),
		(x"00",x"CD",x"4C",x"4F",x"4F",x"4F",x"4E",x"4F",x"4E",x"4E",x"CB",x"CE",x"C8",x"CD",x"CA",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"D3",x"CD",x"C9",x"D0",x"C8",x"CA",x"CC",x"D0",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"01",x"4C",x"CD",x"CC",x"CD",x"CA",x"CD",x"CC",x"01",x"50",x"CB",x"CC",x"CC",x"CA",x"D1",x"C8",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"4D",x"50",x"4E",x"4E",x"4E",x"50",x"4D",x"4E",x"4E",x"CB",x"CE",x"C8",x"CD",x"CA",x"CC",x"00",x"4D",x"CC",x"CB",x"C8",x"CC",x"CF",x"CB",x"01",x"50",x"CB",x"CC",x"CC",x"CA",x"D1",x"C8",x"01",x"4C",x"CD",x"CC",x"CD",x"CA",x"CD",x"CC",x"01",x"50",x"CB",x"CC",x"CC",x"CA",x"D1",x"C8",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"04",x"52",x"CA",x"C9",x"CC",x"CF",x"CD",x"CB",x"00",x"4D",x"D4",x"C0",x"D4",x"CB",x"C8",x"CE",x"00",x"52",x"4D",x"4D",x"50",x"4F",x"51",x"4D",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E"),
		(x"00",x"CD",x"4C",x"4F",x"4F",x"4F",x"4E",x"4F",x"4E",x"4E",x"CB",x"CE",x"C8",x"CD",x"CA",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"C8",x"C8",x"CC",x"CC",x"CB",x"D3",x"CC",x"C7",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"56",x"C5",x"C7",x"C8",x"CC",x"D0",x"CD",x"03",x"4D",x"C6",x"CC",x"CE",x"CD",x"CF",x"CA",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"4D",x"50",x"4E",x"4E",x"4E",x"50",x"4D",x"4E",x"4E",x"CB",x"CE",x"C8",x"CD",x"CA",x"CC",x"00",x"4B",x"D3",x"CE",x"CC",x"CB",x"CA",x"CF",x"03",x"4D",x"C6",x"CC",x"CE",x"CD",x"CF",x"CA",x"00",x"56",x"C5",x"C7",x"C8",x"CC",x"D0",x"CD",x"03",x"4D",x"C6",x"CC",x"CE",x"CD",x"CF",x"CA",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"4F",x"CA",x"CE",x"CB",x"D3",x"CB",x"CF",x"08",x"42",x"CC",x"D0",x"C5",x"CE",x"CC",x"D0",x"02",x"50",x"48",x"4E",x"53",x"51",x"50",x"4F",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E"),
		(x"00",x"CD",x"4C",x"4F",x"4F",x"4F",x"4E",x"4F",x"4E",x"4E",x"CB",x"CE",x"C8",x"CD",x"CA",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"CE",x"C8",x"D0",x"CA",x"CA",x"CF",x"CA",x"D0",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"07",x"49",x"D2",x"CD",x"CD",x"CE",x"CD",x"C9",x"03",x"4F",x"C9",x"CE",x"CD",x"CE",x"D0",x"CA",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"4D",x"50",x"4E",x"4E",x"4E",x"50",x"4D",x"4E",x"4E",x"CB",x"CE",x"C8",x"CD",x"CA",x"CC",x"08",x"47",x"C5",x"D8",x"C9",x"CB",x"CB",x"C9",x"03",x"4F",x"C9",x"CE",x"CD",x"CE",x"D0",x"CA",x"07",x"49",x"D2",x"CD",x"CD",x"CE",x"CD",x"C9",x"03",x"4F",x"C9",x"CE",x"CD",x"CE",x"D0",x"CA",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"54",x"CB",x"C7",x"CE",x"C5",x"CD",x"CC",x"00",x"56",x"CB",x"CE",x"CD",x"C9",x"CC",x"C5",x"01",x"52",x"4D",x"4F",x"50",x"53",x"50",x"4D",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E"),
		(x"00",x"CD",x"4C",x"4F",x"4F",x"4F",x"4E",x"4F",x"4E",x"4E",x"CB",x"CE",x"C8",x"CD",x"CA",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"D0",x"D5",x"C7",x"C9",x"CB",x"D2",x"C8",x"CF",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"4A",x"CB",x"CB",x"CA",x"D1",x"C9",x"C7",x"00",x"4A",x"CD",x"D1",x"C6",x"C7",x"C5",x"D2",x"00",x"4D",x"50",x"4E",x"4E",x"4E",x"50",x"4D",x"4E",x"4E",x"CB",x"CE",x"C8",x"CD",x"CA",x"CC",x"02",x"51",x"CB",x"CF",x"CF",x"C3",x"D1",x"C7",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"4A",x"CB",x"CB",x"CA",x"D1",x"C9",x"C7",x"00",x"4A",x"CD",x"D1",x"C6",x"C7",x"C5",x"D2",x"00",x"4A",x"CB",x"CB",x"CA",x"D1",x"C9",x"C7",x"00",x"4A",x"CD",x"D1",x"C6",x"C7",x"C5",x"D2",x"00",x"4A",x"50",x"50",x"4C",x"4D",x"4C",x"47",x"4D",x"4D",x"51",x"50",x"4C",x"4A",x"4F",x"4E"),
		(x"00",x"CD",x"4C",x"4F",x"4F",x"4F",x"4E",x"4F",x"4E",x"4E",x"CB",x"CE",x"C8",x"CD",x"CA",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"00",x"CF",x"CB",x"CA",x"CB",x"CB",x"C4",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"03",x"51",x"C7",x"CF",x"C7",x"C9",x"D2",x"C8",x"CD",x"C7",x"CC",x"C9",x"C8",x"CF",x"CA",x"CC",x"00",x"4D",x"50",x"4E",x"4E",x"4E",x"50",x"4D",x"4E",x"4E",x"CB",x"CE",x"C8",x"CD",x"CA",x"CC",x"0A",x"CC",x"CB",x"C7",x"D2",x"C5",x"C9",x"CF",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"03",x"51",x"C7",x"CF",x"C7",x"C9",x"D2",x"C8",x"CD",x"C7",x"CC",x"C9",x"C8",x"CF",x"CA",x"CC",x"03",x"51",x"C7",x"CF",x"C7",x"C9",x"D2",x"C8",x"CD",x"C7",x"CC",x"C9",x"C8",x"CF",x"CA",x"CC",x"03",x"58",x"C7",x"C8",x"D1",x"D0",x"CA",x"CD",x"4C",x"4E",x"54",x"51",x"4A",x"4C",x"4F",x"4D"),
		(x"00",x"CD",x"4C",x"4F",x"4F",x"4F",x"4E",x"4F",x"4E",x"4E",x"CB",x"CE",x"C8",x"CD",x"CA",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"0A",x"CA",x"D0",x"CD",x"C6",x"CC",x"D1",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"02",x"47",x"CC",x"CE",x"CD",x"CD",x"CD",x"CC",x"D3",x"CE",x"CA",x"CB",x"D2",x"CA",x"C4",x"D0",x"00",x"4D",x"50",x"4E",x"4E",x"4E",x"50",x"4D",x"4E",x"4E",x"CB",x"CE",x"C8",x"CD",x"CA",x"CC",x"00",x"C8",x"CC",x"CD",x"CA",x"CB",x"CD",x"CD",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"02",x"47",x"CC",x"CE",x"CD",x"CD",x"CD",x"CC",x"D3",x"CE",x"CA",x"CB",x"D2",x"CA",x"C4",x"D0",x"02",x"47",x"CC",x"CE",x"CD",x"CD",x"CD",x"CC",x"D3",x"CE",x"CA",x"CB",x"D2",x"CA",x"C4",x"D0",x"04",x"4B",x"D9",x"CA",x"CD",x"CC",x"CA",x"CE",x"51",x"4C",x"50",x"52",x"4C",x"4D",x"4E",x"4E"),
		(x"00",x"CD",x"4C",x"4F",x"4F",x"4F",x"4E",x"4F",x"4E",x"4E",x"CB",x"CE",x"C8",x"CD",x"CA",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"01",x"03",x"CB",x"CD",x"D3",x"C6",x"CA",x"CA",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"04",x"57",x"C5",x"CB",x"CD",x"C9",x"D3",x"C6",x"C3",x"CD",x"CD",x"CA",x"CA",x"D3",x"C4",x"D5",x"00",x"4D",x"50",x"4E",x"4E",x"4E",x"50",x"4D",x"4E",x"4E",x"CB",x"CE",x"C8",x"CD",x"CA",x"CC",x"01",x"D0",x"C7",x"CC",x"CC",x"CA",x"D0",x"D1",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"04",x"57",x"C5",x"CB",x"CD",x"C9",x"D3",x"C6",x"C3",x"CD",x"CD",x"CA",x"CA",x"D3",x"C4",x"D5",x"04",x"57",x"C5",x"CB",x"CD",x"C9",x"D3",x"C6",x"C3",x"CD",x"CD",x"CA",x"CA",x"D3",x"C4",x"D5",x"00",x"48",x"C3",x"C6",x"C7",x"CB",x"D3",x"CE",x"52",x"49",x"48",x"53",x"50",x"4F",x"4D",x"50"),
		(x"00",x"CD",x"4C",x"4F",x"4F",x"4F",x"4E",x"4F",x"4E",x"4E",x"CB",x"CE",x"C8",x"CD",x"CA",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"02",x"06",x"D0",x"C5",x"CF",x"C7",x"CC",x"CA",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"01",x"4F",x"4E",x"D0",x"C6",x"CA",x"CB",x"D0",x"D0",x"CD",x"C4",x"CF",x"D0",x"C5",x"CF",x"00",x"00",x"4D",x"50",x"4E",x"4E",x"4E",x"50",x"4D",x"4E",x"4E",x"CB",x"CE",x"C8",x"CD",x"CA",x"CC",x"02",x"CA",x"CD",x"C4",x"D2",x"C6",x"CD",x"00",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"01",x"4F",x"4E",x"D0",x"C6",x"CA",x"CB",x"D0",x"D0",x"CD",x"C4",x"CF",x"D0",x"C5",x"CF",x"00",x"01",x"4F",x"4E",x"D0",x"C6",x"CA",x"CB",x"D0",x"D0",x"CD",x"C4",x"CF",x"D0",x"C5",x"CF",x"00",x"00",x"55",x"C7",x"D0",x"CC",x"C9",x"CB",x"C9",x"50",x"5D",x"50",x"53",x"4C",x"4D",x"50",x"52"),
		(x"00",x"CD",x"4C",x"4F",x"4F",x"4F",x"4E",x"4F",x"4E",x"4E",x"CB",x"CE",x"C8",x"CD",x"CA",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"56",x"C0",x"C8",x"D2",x"CD",x"CB",x"CD",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"4D",x"51",x"CA",x"CC",x"CB",x"CD",x"CC",x"C8",x"C5",x"CF",x"D1",x"D0",x"CB",x"CA",x"03",x"00",x"4D",x"50",x"4E",x"4E",x"4E",x"50",x"4D",x"4E",x"4E",x"CB",x"CE",x"C8",x"CD",x"CA",x"CC",x"01",x"D0",x"C9",x"CE",x"D0",x"C6",x"DB",x"00",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"4D",x"51",x"CA",x"CC",x"CB",x"CD",x"CC",x"C8",x"C5",x"CF",x"D1",x"D0",x"CB",x"CA",x"03",x"00",x"4D",x"51",x"CA",x"CC",x"CB",x"CD",x"CC",x"C8",x"C5",x"CF",x"D1",x"D0",x"CB",x"CA",x"03",x"03",x"58",x"D0",x"C9",x"D1",x"CD",x"CB",x"D0",x"00",x"40",x"49",x"54",x"52",x"52",x"53",x"47"),
		(x"00",x"CD",x"4C",x"4F",x"4F",x"4F",x"4E",x"4F",x"4E",x"4E",x"CB",x"CE",x"C8",x"CD",x"CA",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"01",x"56",x"CE",x"C6",x"C7",x"C6",x"CB",x"CF",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"56",x"47",x"00",x"C9",x"CB",x"CC",x"CA",x"D6",x"C9",x"C5",x"CB",x"CB",x"CD",x"00",x"00",x"00",x"4D",x"50",x"4E",x"4E",x"4E",x"50",x"4D",x"4E",x"4E",x"CB",x"CE",x"C8",x"CD",x"CA",x"CC",x"06",x"C7",x"CB",x"CA",x"D0",x"D1",x"00",x"02",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"56",x"47",x"00",x"C9",x"CB",x"CC",x"CA",x"D6",x"C9",x"C5",x"CB",x"CB",x"CD",x"00",x"00",x"00",x"56",x"47",x"00",x"C9",x"CB",x"CC",x"CA",x"D6",x"C9",x"C5",x"CB",x"CB",x"CD",x"00",x"00",x"00",x"4D",x"CC",x"C5",x"CF",x"CD",x"C8",x"C7",x"02",x"58",x"4D",x"4F",x"4A",x"49",x"56",x"50"),
		(x"00",x"CD",x"4C",x"4F",x"4F",x"4F",x"4E",x"4F",x"4E",x"4E",x"CB",x"CE",x"C8",x"CD",x"CA",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"03",x"47",x"CB",x"C8",x"D1",x"CF",x"CA",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"01",x"4C",x"4D",x"02",x"CE",x"C9",x"D3",x"CB",x"C8",x"D3",x"C7",x"CD",x"C8",x"C9",x"02",x"00",x"00",x"4D",x"50",x"4E",x"4E",x"4E",x"50",x"4D",x"4E",x"4E",x"CB",x"CE",x"C8",x"CD",x"CA",x"CC",x"01",x"C2",x"D4",x"CA",x"CA",x"CF",x"00",x"07",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"00",x"50",x"CC",x"CB",x"CB",x"CE",x"C9",x"CC",x"01",x"4C",x"4D",x"02",x"CE",x"C9",x"D3",x"CB",x"C8",x"D3",x"C7",x"CD",x"C8",x"C9",x"02",x"00",x"01",x"4C",x"4D",x"02",x"CE",x"C9",x"D3",x"CB",x"C8",x"D3",x"C7",x"CD",x"C8",x"C9",x"02",x"00",x"00",x"52",x"C9",x"CE",x"C9",x"C9",x"D2",x"CE",x"00",x"57",x"46",x"55",x"56",x"47",x"52",x"4D"),
		(x"02",x"CD",x"48",x"4C",x"50",x"4D",x"4F",x"4C",x"52",x"51",x"C4",x"CD",x"D8",x"CF",x"C4",x"C9",x"00",x"53",x"CB",x"CF",x"C4",x"CD",x"D4",x"C4",x"00",x"53",x"CB",x"CF",x"C4",x"CD",x"D4",x"C4",x"00",x"53",x"CB",x"CF",x"C4",x"CD",x"D4",x"C4",x"00",x"53",x"CB",x"CF",x"C4",x"CD",x"D4",x"C4",x"00",x"53",x"CB",x"CF",x"C4",x"CD",x"D4",x"C4",x"00",x"53",x"CB",x"CF",x"C4",x"CD",x"D4",x"C4",x"00",x"53",x"CB",x"CF",x"C4",x"CD",x"D4",x"C4",x"04",x"47",x"53",x"46",x"02",x"CB",x"C9",x"CD",x"CA",x"CD",x"D2",x"BF",x"C6",x"06",x"03",x"00",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"52",x"51",x"C4",x"CD",x"D8",x"CF",x"C4",x"C9",x"00",x"CC",x"C1",x"D2",x"C5",x"06",x"00",x"00",x"52",x"51",x"C4",x"CD",x"D8",x"CF",x"C4",x"C9",x"00",x"53",x"CB",x"CF",x"C4",x"CD",x"D4",x"C4",x"04",x"47",x"53",x"46",x"02",x"CB",x"C9",x"CD",x"CA",x"CD",x"D2",x"BF",x"C6",x"06",x"03",x"00",x"51",x"56",x"4E",x"55",x"08",x"C9",x"C7",x"CB",x"CA",x"CD",x"D2",x"BF",x"C6",x"06",x"03",x"00",x"52",x"51",x"C4",x"CD",x"D8",x"CF",x"C4",x"C9",x"02",x"4C",x"4B",x"4D",x"4D",x"4F",x"4F",x"54"),
		(x"09",x"C2",x"54",x"49",x"51",x"4C",x"50",x"53",x"46",x"53",x"52",x"00",x"00",x"01",x"00",x"03",x"00",x"4B",x"4F",x"00",x"00",x"08",x"06",x"00",x"00",x"4B",x"4F",x"00",x"00",x"08",x"06",x"00",x"00",x"4B",x"4F",x"00",x"00",x"08",x"06",x"00",x"00",x"4B",x"4F",x"00",x"00",x"08",x"06",x"00",x"00",x"4B",x"4F",x"00",x"00",x"08",x"06",x"00",x"00",x"4B",x"4F",x"00",x"00",x"08",x"06",x"00",x"00",x"4B",x"4F",x"00",x"00",x"08",x"06",x"00",x"00",x"4F",x"53",x"54",x"06",x"06",x"05",x"01",x"01",x"04",x"00",x"00",x"00",x"03",x"02",x"00",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"46",x"53",x"52",x"00",x"00",x"01",x"00",x"03",x"06",x"55",x"08",x"07",x"07",x"04",x"00",x"06",x"46",x"53",x"52",x"00",x"00",x"01",x"00",x"03",x"00",x"4B",x"4F",x"00",x"00",x"08",x"06",x"00",x"00",x"4F",x"53",x"54",x"06",x"06",x"05",x"01",x"01",x"04",x"00",x"00",x"00",x"03",x"02",x"00",x"4C",x"47",x"4B",x"47",x"00",x"05",x"08",x"04",x"01",x"04",x"00",x"00",x"00",x"03",x"02",x"00",x"46",x"53",x"52",x"00",x"00",x"01",x"00",x"03",x"00",x"4C",x"55",x"4F",x"4E",x"4A",x"4F",x"4A"),
		(x"00",x"CD",x"4E",x"53",x"4F",x"4F",x"56",x"49",x"4B",x"53",x"4C",x"00",x"01",x"00",x"00",x"05",x"08",x"4B",x"57",x"07",x"02",x"00",x"06",x"02",x"08",x"4B",x"57",x"07",x"02",x"00",x"06",x"02",x"08",x"4B",x"57",x"07",x"02",x"00",x"06",x"02",x"08",x"4B",x"57",x"07",x"02",x"00",x"06",x"02",x"08",x"4B",x"57",x"07",x"02",x"00",x"06",x"02",x"08",x"4B",x"57",x"07",x"02",x"00",x"06",x"02",x"08",x"4B",x"57",x"07",x"02",x"00",x"06",x"02",x"03",x"57",x"4D",x"44",x"51",x"00",x"00",x"06",x"00",x"0B",x"03",x"06",x"02",x"00",x"00",x"4F",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4B",x"53",x"4C",x"00",x"01",x"00",x"00",x"05",x"00",x"49",x"08",x"0B",x"00",x"00",x"00",x"4F",x"4B",x"53",x"4C",x"00",x"01",x"00",x"00",x"05",x"08",x"4B",x"57",x"07",x"02",x"00",x"06",x"02",x"03",x"57",x"4D",x"44",x"51",x"00",x"00",x"06",x"00",x"0B",x"03",x"06",x"02",x"00",x"00",x"4F",x"50",x"4C",x"50",x"55",x"4A",x"00",x"00",x"10",x"00",x"0B",x"03",x"06",x"02",x"00",x"00",x"4F",x"4B",x"53",x"4C",x"00",x"01",x"00",x"00",x"05",x"00",x"52",x"51",x"4E",x"54",x"4E",x"49",x"57"),
		(x"00",x"C5",x"53",x"59",x"4C",x"46",x"4B",x"53",x"4C",x"4F",x"57",x"00",x"00",x"01",x"00",x"04",x"00",x"4B",x"4A",x"00",x"01",x"00",x"05",x"03",x"00",x"4B",x"4A",x"00",x"01",x"00",x"05",x"03",x"00",x"4B",x"4A",x"00",x"01",x"00",x"05",x"03",x"00",x"4B",x"4A",x"00",x"01",x"00",x"05",x"03",x"00",x"4B",x"4A",x"00",x"01",x"00",x"05",x"03",x"00",x"4B",x"4A",x"00",x"01",x"00",x"05",x"03",x"00",x"4B",x"4A",x"00",x"01",x"00",x"05",x"03",x"00",x"43",x"51",x"4C",x"54",x"00",x"05",x"02",x"03",x"00",x"00",x"06",x"00",x"04",x"04",x"4D",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4C",x"4F",x"57",x"00",x"00",x"01",x"00",x"04",x"06",x"4D",x"01",x"00",x"00",x"01",x"07",x"56",x"4C",x"4F",x"57",x"00",x"00",x"01",x"00",x"04",x"00",x"4B",x"4A",x"00",x"01",x"00",x"05",x"03",x"00",x"43",x"51",x"4C",x"54",x"00",x"05",x"02",x"03",x"00",x"00",x"06",x"00",x"04",x"04",x"4D",x"54",x"4E",x"4F",x"4E",x"4B",x"00",x"00",x"00",x"03",x"00",x"00",x"06",x"00",x"04",x"04",x"4D",x"4C",x"4F",x"57",x"00",x"00",x"01",x"00",x"04",x"00",x"4A",x"4E",x"50",x"52",x"51",x"47",x"44"),
		(x"01",x"CE",x"4E",x"49",x"CF",x"C1",x"54",x"4C",x"50",x"5A",x"4A",x"04",x"01",x"00",x"00",x"03",x"00",x"59",x"55",x"00",x"00",x"05",x"04",x"00",x"00",x"59",x"55",x"00",x"00",x"05",x"04",x"00",x"00",x"59",x"55",x"00",x"00",x"05",x"04",x"00",x"00",x"59",x"55",x"00",x"00",x"05",x"04",x"00",x"00",x"59",x"55",x"00",x"00",x"05",x"04",x"00",x"00",x"59",x"55",x"00",x"00",x"05",x"04",x"00",x"00",x"59",x"55",x"00",x"00",x"05",x"04",x"00",x"07",x"52",x"4F",x"4F",x"44",x"58",x"00",x"01",x"03",x"02",x"00",x"00",x"08",x"00",x"4D",x"54",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"50",x"5A",x"4A",x"04",x"01",x"00",x"00",x"03",x"01",x"47",x"00",x"00",x"0A",x"06",x"4A",x"44",x"50",x"5A",x"4A",x"04",x"01",x"00",x"00",x"03",x"00",x"59",x"55",x"00",x"00",x"05",x"04",x"00",x"07",x"52",x"4F",x"4F",x"44",x"58",x"00",x"01",x"03",x"02",x"00",x"00",x"08",x"00",x"4D",x"54",x"49",x"50",x"4F",x"55",x"4C",x"52",x"00",x"03",x"03",x"02",x"00",x"00",x"08",x"00",x"4D",x"54",x"50",x"5A",x"4A",x"04",x"01",x"00",x"00",x"03",x"09",x"40",x"53",x"49",x"CE",x"CC",x"53",x"50"),
		(x"03",x"C7",x"53",x"4D",x"C3",x"D8",x"04",x"4B",x"4B",x"4F",x"45",x"54",x"55",x"4D",x"4E",x"50",x"59",x"49",x"4A",x"49",x"51",x"4B",x"50",x"4A",x"59",x"49",x"4A",x"49",x"51",x"4B",x"50",x"4A",x"59",x"49",x"4A",x"49",x"51",x"4B",x"50",x"4A",x"59",x"49",x"4A",x"49",x"51",x"4B",x"50",x"4A",x"59",x"49",x"4A",x"49",x"51",x"4B",x"50",x"4A",x"59",x"49",x"4A",x"49",x"51",x"4B",x"50",x"4A",x"59",x"49",x"4A",x"49",x"51",x"4B",x"50",x"4A",x"55",x"4A",x"4F",x"58",x"53",x"49",x"53",x"4A",x"53",x"53",x"4C",x"4E",x"4D",x"54",x"43",x"4D",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4B",x"4F",x"45",x"54",x"55",x"4D",x"4E",x"50",x"4C",x"55",x"52",x"52",x"50",x"4A",x"5A",x"4C",x"4B",x"4F",x"45",x"54",x"55",x"4D",x"4E",x"50",x"59",x"49",x"4A",x"49",x"51",x"4B",x"50",x"4A",x"55",x"4A",x"4F",x"58",x"53",x"49",x"53",x"4A",x"53",x"53",x"4C",x"4E",x"4D",x"54",x"43",x"4D",x"50",x"4C",x"50",x"50",x"4F",x"45",x"54",x"48",x"53",x"53",x"4C",x"4E",x"4D",x"54",x"43",x"4D",x"4B",x"4F",x"45",x"54",x"55",x"4D",x"4E",x"50",x"52",x"55",x"4B",x"4A",x"D0",x"D3",x"00",x"51"),
		(x"01",x"C5",x"56",x"4D",x"4D",x"00",x"05",x"49",x"51",x"4C",x"49",x"57",x"4C",x"52",x"57",x"48",x"4E",x"4C",x"54",x"4D",x"50",x"55",x"4F",x"47",x"4E",x"4C",x"54",x"4D",x"50",x"55",x"4F",x"47",x"4E",x"4C",x"54",x"4D",x"50",x"55",x"4F",x"47",x"4E",x"4C",x"54",x"4D",x"50",x"55",x"4F",x"47",x"4E",x"4C",x"54",x"4D",x"50",x"55",x"4F",x"47",x"4E",x"4C",x"54",x"4D",x"50",x"55",x"4F",x"47",x"4E",x"4C",x"54",x"4D",x"50",x"55",x"4F",x"47",x"4F",x"48",x"55",x"4A",x"58",x"4B",x"4C",x"51",x"4E",x"4C",x"53",x"53",x"4C",x"53",x"50",x"47",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"51",x"4C",x"49",x"57",x"4C",x"52",x"57",x"48",x"53",x"45",x"52",x"48",x"4D",x"4E",x"44",x"4E",x"51",x"4C",x"49",x"57",x"4C",x"52",x"57",x"48",x"4E",x"4C",x"54",x"4D",x"50",x"55",x"4F",x"47",x"4F",x"48",x"55",x"4A",x"58",x"4B",x"4C",x"51",x"4E",x"4C",x"53",x"53",x"4C",x"53",x"50",x"47",x"52",x"4F",x"4D",x"4E",x"52",x"4A",x"4F",x"57",x"4E",x"4C",x"53",x"53",x"4C",x"53",x"50",x"47",x"51",x"4C",x"49",x"57",x"4C",x"52",x"57",x"48",x"45",x"50",x"4F",x"45",x"53",x"00",x"03",x"4F"),
		(x"02",x"D1",x"4A",x"50",x"52",x"4F",x"4B",x"56",x"4F",x"4D",x"57",x"43",x"4F",x"53",x"46",x"51",x"50",x"49",x"54",x"52",x"4B",x"4C",x"4B",x"57",x"50",x"49",x"54",x"52",x"4B",x"4C",x"4B",x"57",x"50",x"49",x"54",x"52",x"4B",x"4C",x"4B",x"57",x"50",x"49",x"54",x"52",x"4B",x"4C",x"4B",x"57",x"50",x"49",x"54",x"52",x"4B",x"4C",x"4B",x"57",x"50",x"49",x"54",x"52",x"4B",x"4C",x"4B",x"57",x"50",x"49",x"54",x"52",x"4B",x"4C",x"4B",x"57",x"4D",x"52",x"4C",x"4F",x"47",x"53",x"50",x"4E",x"4D",x"4E",x"4D",x"53",x"4C",x"48",x"4B",x"58",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4E",x"4F",x"4D",x"57",x"43",x"4F",x"53",x"46",x"51",x"4B",x"4E",x"4E",x"50",x"56",x"47",x"59",x"50",x"4F",x"4D",x"57",x"43",x"4F",x"53",x"46",x"51",x"50",x"49",x"54",x"52",x"4B",x"4C",x"4B",x"57",x"4D",x"52",x"4C",x"4F",x"47",x"53",x"50",x"4E",x"4D",x"4E",x"4D",x"53",x"4C",x"48",x"4B",x"58",x"4C",x"4B",x"4F",x"54",x"4C",x"4E",x"4E",x"50",x"4D",x"4E",x"4D",x"53",x"4C",x"48",x"4B",x"58",x"4F",x"4D",x"57",x"43",x"4F",x"53",x"46",x"51",x"51",x"4D",x"51",x"53",x"4B",x"4C",x"4D",x"4F")
	
	);
	
	constant titulo_B : ROM :=
	(
		
		(x"EA",x"DE",x"D5",x"D7",x"DD",x"DD",x"DA",x"DA",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"DC",x"D8",x"D6",x"E9",x"E0",x"D4",x"D5",x"E3",x"DB"),
		(x"DD",x"C8",x"C7",x"CF",x"CC",x"C2",x"D4",x"BB",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C0",x"BC",x"B9",x"D5",x"C9",x"C8",x"BD",x"C1"),
		(x"D1",x"CE",x"00",x"00",x"09",x"00",x"0B",x"06",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"10",x"00",x"08",x"00",x"03",x"06",x"09",x"00"),
		(x"D1",x"CF",x"00",x"00",x"06",x"03",x"00",x"00",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"05",x"16",x"00",x"03",x"06",x"01",x"00",x"07"),
		(x"E2",x"CB",x"05",x"0C",x"C6",x"C5",x"00",x"05",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"06",x"00",x"00",x"BE",x"BD",x"00",x"05"),
		(x"E3",x"BE",x"00",x"02",x"C4",x"D8",x"04",x"03",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"00",x"06",x"06",x"05",x"C0",x"E5",x"06",x"00"),
		(x"D5",x"D6",x"11",x"00",x"00",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"07",x"00",x"05",x"00",x"00",x"00",x"00",x"00"),
		(x"D9",x"BD",x"08",x"00",x"07",x"06",x"00",x"16",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"00",x"01",x"00",x"00",x"0C",x"00",x"00",x"0A"),
		(x"DC",x"C1",x"03",x"02",x"00",x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"07",x"05",x"00",x"00",x"00",x"17",x"00",x"00",x"00",x"00",x"04",x"00",x"1C",x"09",x"00",x"00",x"03",x"00",x"06",x"00",x"0D",x"00",x"00",x"00",x"03",x"00",x"06",x"00",x"0D",x"00",x"00",x"00",x"03",x"00",x"00",x"00",x"00",x"17",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"07",x"05",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"06",x"00",x"0D",x"00",x"00",x"00",x"03",x"00",x"00",x"00",x"00",x"17",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"DC",x"C1",x"03",x"02",x"00",x"02",x"00",x"00",x"00",x"12",x"0D",x"00",x"0D",x"D0",x"C7",x"BA",x"DE",x"BE",x"BC",x"CD",x"C6",x"00",x"00",x"06",x"00",x"08",x"AF",x"B3",x"C3",x"C2",x"CA",x"CC",x"00",x"15",x"B8",x"C8",x"D1",x"CC",x"D1",x"C9",x"00",x"15",x"B8",x"C8",x"D1",x"CC",x"D1",x"C9",x"DE",x"BE",x"BC",x"CD",x"C6",x"00",x"00",x"06",x"00",x"12",x"0D",x"00",x"0D",x"D0",x"C7",x"BA",x"C8",x"C8",x"C8",x"C8",x"C8",x"C8",x"C8",x"C8",x"00",x"15",x"B8",x"C8",x"D1",x"CC",x"D1",x"C9",x"DE",x"BE",x"BC",x"CD",x"C6",x"00",x"00",x"06",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"DC",x"C1",x"03",x"02",x"00",x"02",x"00",x"00",x"00",x"00",x"07",x"08",x"C2",x"C8",x"BC",x"CE",x"C4",x"BB",x"C7",x"B1",x"C6",x"CA",x"00",x"05",x"00",x"00",x"CB",x"C6",x"CE",x"C5",x"C5",x"BF",x"04",x"00",x"C8",x"C9",x"C8",x"C0",x"BC",x"B5",x"04",x"00",x"C8",x"C9",x"C8",x"C0",x"BC",x"B5",x"C4",x"BB",x"C7",x"B1",x"C6",x"CA",x"00",x"05",x"00",x"00",x"07",x"08",x"C2",x"C8",x"BC",x"CE",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"04",x"00",x"C8",x"C9",x"C8",x"C0",x"BC",x"B5",x"C4",x"BB",x"C7",x"B1",x"C6",x"CA",x"00",x"05",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"DC",x"C1",x"03",x"02",x"00",x"02",x"00",x"00",x"0B",x"06",x"09",x"00",x"BA",x"B0",x"C9",x"B7",x"CF",x"BD",x"C5",x"D2",x"C3",x"CC",x"03",x"07",x"08",x"0A",x"C5",x"CC",x"CD",x"C2",x"C4",x"B5",x"10",x"00",x"C9",x"CB",x"C4",x"C1",x"C3",x"CF",x"10",x"00",x"C9",x"CB",x"C4",x"C1",x"C3",x"CF",x"CF",x"BD",x"C5",x"D2",x"C3",x"CC",x"03",x"07",x"0B",x"06",x"09",x"00",x"BA",x"B0",x"C9",x"B7",x"C4",x"C4",x"C4",x"C4",x"C4",x"C4",x"C4",x"C4",x"10",x"00",x"C9",x"CB",x"C4",x"C1",x"C3",x"CF",x"CF",x"BD",x"C5",x"D2",x"C3",x"CC",x"03",x"07",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"DC",x"C1",x"03",x"02",x"00",x"02",x"00",x"00",x"00",x"07",x"00",x"C2",x"D1",x"D0",x"BC",x"C7",x"B6",x"D0",x"C3",x"C2",x"D4",x"B8",x"CA",x"05",x"00",x"0E",x"BC",x"CA",x"CC",x"C4",x"CD",x"C6",x"00",x"00",x"BA",x"C4",x"C2",x"CD",x"C5",x"CD",x"00",x"00",x"BA",x"C4",x"C2",x"CD",x"C5",x"CD",x"B6",x"D0",x"C3",x"C2",x"D4",x"B8",x"CA",x"05",x"00",x"07",x"00",x"C2",x"D1",x"D0",x"BC",x"C7",x"C7",x"C7",x"C7",x"C7",x"C7",x"C7",x"C7",x"C7",x"00",x"00",x"BA",x"C4",x"C2",x"CD",x"C5",x"CD",x"B6",x"D0",x"C3",x"C2",x"D4",x"B8",x"CA",x"05",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"DC",x"C1",x"03",x"02",x"00",x"02",x"00",x"00",x"0C",x"04",x"00",x"D0",x"CF",x"B9",x"C6",x"E1",x"C5",x"D8",x"CC",x"BA",x"B6",x"CE",x"C5",x"00",x"00",x"00",x"B4",x"B1",x"C1",x"BE",x"C7",x"CB",x"00",x"02",x"D2",x"D0",x"B8",x"C2",x"BC",x"C8",x"00",x"02",x"D2",x"D0",x"B8",x"C2",x"BC",x"C8",x"C5",x"D8",x"CC",x"BA",x"B6",x"CE",x"C5",x"00",x"0C",x"04",x"00",x"D0",x"CF",x"B9",x"C6",x"E1",x"C7",x"C7",x"C7",x"C7",x"C7",x"C7",x"C7",x"C7",x"00",x"02",x"D2",x"D0",x"B8",x"C2",x"BC",x"C8",x"C5",x"D8",x"CC",x"BA",x"B6",x"CE",x"C5",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"DC",x"C1",x"03",x"02",x"00",x"02",x"00",x"00",x"00",x"00",x"B7",x"C2",x"C9",x"BD",x"D1",x"AB",x"B8",x"BA",x"CA",x"D8",x"BB",x"CA",x"BB",x"D0",x"0A",x"08",x"C2",x"C0",x"CD",x"C4",x"C3",x"BC",x"0B",x"0C",x"C5",x"BC",x"B2",x"CB",x"CC",x"D1",x"0B",x"0C",x"C5",x"BC",x"B2",x"CB",x"CC",x"D1",x"B8",x"BA",x"CA",x"D8",x"BB",x"CA",x"BB",x"D0",x"00",x"00",x"B7",x"C2",x"C9",x"BD",x"D1",x"AB",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"C1",x"0B",x"0C",x"C5",x"BC",x"B2",x"CB",x"CC",x"D1",x"B8",x"BA",x"CA",x"D8",x"BB",x"CA",x"BB",x"D0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"DC",x"C1",x"03",x"02",x"00",x"02",x"00",x"00",x"03",x"00",x"D1",x"C7",x"B5",x"D0",x"C3",x"C1",x"C9",x"CE",x"C5",x"BB",x"D6",x"C6",x"B7",x"CF",x"00",x"05",x"BF",x"CE",x"CC",x"C3",x"CA",x"BC",x"00",x"00",x"C8",x"D0",x"C8",x"CF",x"BF",x"BA",x"00",x"00",x"C8",x"D0",x"C8",x"CF",x"BF",x"BA",x"C9",x"CE",x"C5",x"BB",x"D6",x"C6",x"B7",x"CF",x"03",x"00",x"D1",x"C7",x"B5",x"D0",x"C3",x"C1",x"C8",x"C8",x"C8",x"C8",x"C8",x"C8",x"C8",x"C8",x"00",x"00",x"C8",x"D0",x"C8",x"CF",x"BF",x"BA",x"C9",x"CE",x"C5",x"BB",x"D6",x"C6",x"B7",x"CF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"DC",x"C1",x"03",x"02",x"00",x"02",x"00",x"00",x"04",x"00",x"CF",x"D6",x"B7",x"D2",x"CC",x"BA",x"C8",x"C4",x"BE",x"BF",x"C4",x"C8",x"CB",x"CC",x"00",x"00",x"C8",x"C8",x"C7",x"BF",x"C4",x"C5",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"D2",x"C1",x"C3",x"CA",x"C7",x"C3",x"BE",x"CA",x"2D",x"00",x"BF",x"C3",x"C7",x"C6",x"C6",x"C8",x"CD",x"C6",x"BF",x"C0",x"CB",x"CF",x"C2",x"B7",x"0A",x"00",x"BC",x"C8",x"C1",x"CB",x"B9",x"C6",x"C9",x"BC",x"C0",x"C6",x"CE",x"C5",x"C2",x"C4",x"2C",x"00",x"00",x"03",x"00",x"00",x"02",x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"DC",x"C1",x"03",x"02",x"00",x"02",x"00",x"00",x"04",x"00",x"D7",x"B4",x"C8",x"B1",x"D5",x"C4",x"C1",x"06",x"13",x"07",x"00",x"00",x"02",x"00",x"10",x"07",x"BE",x"C2",x"CB",x"C5",x"C9",x"C8",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"00",x"CA",x"BA",x"C1",x"C9",x"C6",x"C0",x"C3",x"00",x"00",x"CD",x"C4",x"C4",x"C7",x"C7",x"C1",x"02",x"00",x"00",x"05",x"09",x"04",x"00",x"0B",x"09",x"00",x"BA",x"C7",x"C3",x"C9",x"B9",x"C9",x"00",x"CB",x"B9",x"CC",x"CB",x"C4",x"C4",x"C1",x"00",x"00",x"06",x"02",x"00",x"01",x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"DC",x"C1",x"03",x"02",x"00",x"02",x"00",x"00",x"00",x"0C",x"BF",x"B3",x"C9",x"B8",x"CC",x"C0",x"BD",x"D1",x"09",x"00",x"00",x"12",x"0B",x"00",x"00",x"19",x"C8",x"B9",x"C4",x"C8",x"BC",x"BC",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"00",x"C7",x"C3",x"CB",x"C4",x"BC",x"C3",x"CD",x"00",x"07",x"D6",x"C3",x"C5",x"C1",x"C4",x"C7",x"09",x"BB",x"B7",x"CD",x"BB",x"B0",x"D2",x"15",x"00",x"08",x"C1",x"C8",x"C2",x"C5",x"BF",x"CA",x"07",x"C6",x"CE",x"C6",x"C4",x"B7",x"BF",x"CA",x"00",x"09",x"0F",x"00",x"00",x"00",x"00",x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"DC",x"C1",x"03",x"02",x"00",x"02",x"00",x"00",x"06",x"0A",x"09",x"CA",x"BA",x"C8",x"BF",x"C1",x"CB",x"BF",x"B8",x"C6",x"00",x"05",x"07",x"00",x"00",x"00",x"BE",x"C4",x"C1",x"D3",x"CB",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"00",x"C6",x"C1",x"C9",x"CB",x"C4",x"C8",x"CC",x"05",x"0B",x"CD",x"C3",x"CD",x"C0",x"C5",x"C8",x"00",x"CB",x"C9",x"D1",x"D0",x"BA",x"B7",x"00",x"00",x"12",x"C8",x"C7",x"C1",x"C2",x"C4",x"CB",x"05",x"CF",x"BB",x"C5",x"C8",x"C6",x"C6",x"C9",x"04",x"0C",x"06",x"01",x"06",x"00",x"00",x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"DC",x"C1",x"03",x"02",x"00",x"02",x"00",x"00",x"15",x"00",x"00",x"C0",x"CF",x"BB",x"D1",x"CA",x"BF",x"C4",x"CB",x"C9",x"C7",x"D7",x"00",x"00",x"00",x"00",x"D9",x"CF",x"BE",x"CA",x"B3",x"BC",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"03",x"C6",x"C9",x"BA",x"C7",x"C3",x"C8",x"00",x"00",x"02",x"C8",x"BF",x"C4",x"C4",x"CE",x"C4",x"00",x"C9",x"C1",x"BD",x"C9",x"D7",x"D4",x"00",x"00",x"00",x"BD",x"C8",x"C8",x"C2",x"C4",x"C9",x"0A",x"C4",x"C2",x"C5",x"C0",x"C6",x"C8",x"02",x"00",x"04",x"02",x"00",x"00",x"00",x"0B",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"DC",x"C1",x"03",x"02",x"00",x"02",x"00",x"00",x"00",x"00",x"00",x"0C",x"CF",x"CC",x"B9",x"BE",x"BF",x"C7",x"D0",x"BC",x"BB",x"CA",x"B3",x"1B",x"18",x"00",x"C1",x"D7",x"C7",x"C8",x"C7",x"CF",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"04",x"CC",x"BE",x"CB",x"C9",x"C3",x"D1",x"00",x"00",x"01",x"C6",x"BC",x"BF",x"C4",x"D3",x"C4",x"00",x"CF",x"C6",x"C2",x"CD",x"B7",x"B0",x"10",x"1F",x"18",x"C1",x"C7",x"C6",x"B9",x"C1",x"D1",x"00",x"C7",x"C0",x"BB",x"CD",x"C9",x"00",x"00",x"00",x"03",x"00",x"00",x"00",x"00",x"0F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"DC",x"C1",x"03",x"02",x"00",x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"06",x"C8",x"C4",x"BC",x"D1",x"B9",x"C1",x"C2",x"CA",x"A9",x"0A",x"07",x"00",x"BF",x"C7",x"C8",x"C2",x"C3",x"C0",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"C9",x"C0",x"C5",x"C8",x"C9",x"00",x"03",x"00",x"00",x"C1",x"BF",x"CC",x"C9",x"C8",x"BD",x"00",x"C1",x"B8",x"BA",x"C5",x"C6",x"C9",x"00",x"03",x"00",x"B9",x"CC",x"D0",x"C1",x"BF",x"C5",x"03",x"CC",x"BF",x"C3",x"CC",x"BF",x"CB",x"00",x"00",x"00",x"00",x"00",x"06",x"03",x"03",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"DC",x"C1",x"03",x"02",x"00",x"02",x"00",x"00",x"15",x"05",x"05",x"00",x"01",x"02",x"05",x"00",x"C9",x"C5",x"C9",x"C5",x"C8",x"C8",x"CA",x"B8",x"04",x"05",x"B4",x"BC",x"CB",x"C7",x"D5",x"C0",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"05",x"C7",x"BE",x"C4",x"CD",x"C6",x"00",x"05",x"01",x"04",x"CB",x"BD",x"CB",x"C7",x"C3",x"BF",x"09",x"CD",x"C9",x"CE",x"C9",x"B9",x"C1",x"0E",x"00",x"00",x"BE",x"C7",x"C8",x"C2",x"C4",x"C6",x"03",x"C6",x"C3",x"CE",x"C4",x"C4",x"C4",x"CB",x"02",x"07",x"05",x"00",x"04",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"DC",x"C1",x"03",x"02",x"00",x"02",x"00",x"00",x"01",x"02",x"01",x"09",x"00",x"0B",x"04",x"00",x"00",x"00",x"C5",x"C8",x"C7",x"C7",x"CC",x"BC",x"00",x"00",x"D0",x"C2",x"C4",x"C7",x"BA",x"C9",x"00",x"18",x"C7",x"D1",x"B4",x"CE",x"C3",x"C5",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"00",x"D7",x"B1",x"D2",x"BC",x"00",x"02",x"03",x"00",x"05",x"C8",x"C2",x"C4",x"C5",x"C1",x"C7",x"00",x"1A",x"00",x"00",x"00",x"07",x"07",x"00",x"00",x"07",x"C4",x"C7",x"C9",x"BF",x"CD",x"C6",x"15",x"98",x"D4",x"C4",x"C9",x"C7",x"C0",x"BF",x"00",x"00",x"00",x"01",x"03",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"DC",x"C1",x"03",x"02",x"00",x"02",x"00",x"00",x"07",x"00",x"BB",x"AF",x"C4",x"CA",x"C6",x"D1",x"C9",x"D1",x"C8",x"C4",x"C8",x"C7",x"B9",x"C8",x"04",x"00",x"C8",x"CD",x"C7",x"BF",x"BD",x"C9",x"C4",x"AA",x"C5",x"C3",x"B7",x"D3",x"CE",x"B9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"00",x"00",x"08",x"07",x"02",x"1A",x"00",x"00",x"04",x"0B",x"C2",x"CA",x"C4",x"BF",x"CB",x"C8",x"C6",x"AE",x"CE",x"CE",x"BC",x"D6",x"CB",x"D1",x"00",x"04",x"C7",x"C7",x"C9",x"C2",x"CA",x"C4",x"07",x"10",x"D2",x"BF",x"C4",x"C8",x"C5",x"C5",x"02",x"00",x"00",x"07",x"0D",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"DC",x"C1",x"03",x"02",x"00",x"02",x"00",x"00",x"00",x"01",x"CB",x"D3",x"BB",x"B8",x"B5",x"C0",x"CD",x"C9",x"C1",x"C4",x"C7",x"CA",x"C9",x"CB",x"1B",x"0D",x"C7",x"C6",x"C5",x"C6",x"BD",x"D4",x"C6",x"CA",x"C3",x"BE",x"C4",x"CA",x"CA",x"BC",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"0B",x"00",x"00",x"06",x"00",x"02",x"16",x"00",x"00",x"BC",x"CA",x"CB",x"C6",x"C8",x"C9",x"C4",x"C4",x"CB",x"C4",x"D0",x"C5",x"BA",x"C2",x"03",x"00",x"C1",x"C7",x"C8",x"C5",x"C6",x"C3",x"01",x"00",x"CA",x"C1",x"BF",x"CC",x"C5",x"C7",x"1E",x"14",x"00",x"02",x"02",x"00",x"00",x"0C",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"DC",x"C1",x"03",x"02",x"00",x"02",x"00",x"00",x"00",x"00",x"B2",x"CE",x"CC",x"D0",x"C5",x"C1",x"C1",x"CC",x"CA",x"C6",x"C4",x"BE",x"C7",x"C4",x"00",x"06",x"A8",x"CA",x"C7",x"C4",x"C8",x"C5",x"B8",x"D3",x"C6",x"B9",x"C2",x"CF",x"C0",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"02",x"00",x"09",x"0A",x"00",x"11",x"03",x"0B",x"A3",x"C6",x"CB",x"C1",x"CB",x"C0",x"B5",x"E5",x"B7",x"BC",x"D5",x"BC",x"BD",x"BC",x"0E",x"00",x"B9",x"C6",x"CB",x"CA",x"C1",x"C3",x"00",x"07",x"BD",x"BF",x"BD",x"CD",x"C6",x"C7",x"00",x"00",x"00",x"03",x"05",x"00",x"00",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"DC",x"C1",x"03",x"02",x"00",x"02",x"00",x"00",x"00",x"07",x"0F",x"BD",x"CD",x"B6",x"CF",x"C5",x"CA",x"C5",x"C3",x"C2",x"C3",x"C4",x"C7",x"00",x"00",x"0A",x"07",x"C1",x"C7",x"D3",x"C5",x"B8",x"CC",x"CE",x"BD",x"C0",x"CF",x"C1",x"BE",x"00",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"09",x"00",x"01",x"04",x"08",x"00",x"00",x"00",x"00",x"00",x"1B",x"C7",x"C2",x"C0",x"C1",x"C4",x"BD",x"D0",x"B5",x"CB",x"CB",x"BF",x"CA",x"C9",x"21",x"06",x"C5",x"C5",x"C3",x"CA",x"C1",x"C5",x"00",x"00",x"C8",x"C1",x"C7",x"C8",x"C7",x"C3",x"00",x"0C",x"07",x"02",x"00",x"00",x"00",x"06",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"DC",x"C1",x"03",x"02",x"00",x"02",x"00",x"00",x"00",x"0A",x"09",x"C1",x"C8",x"B7",x"C7",x"C5",x"BB",x"C7",x"C3",x"CA",x"C0",x"BE",x"D3",x"00",x"07",x"03",x"00",x"C4",x"CE",x"C8",x"C7",x"BE",x"C2",x"C5",x"C8",x"C6",x"D2",x"C5",x"BA",x"0D",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"09",x"00",x"00",x"05",x"00",x"0C",x"00",x"08",x"00",x"00",x"0F",x"BE",x"C7",x"C4",x"C2",x"C0",x"C5",x"C7",x"C1",x"CF",x"C8",x"BE",x"CF",x"C6",x"00",x"00",x"C1",x"C7",x"C4",x"D0",x"C2",x"BD",x"05",x"06",x"D0",x"C2",x"C9",x"C5",x"C7",x"BE",x"00",x"04",x"00",x"02",x"00",x"02",x"00",x"05",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"DC",x"C1",x"03",x"02",x"00",x"02",x"00",x"00",x"03",x"00",x"0A",x"00",x"BC",x"BC",x"C6",x"C3",x"BF",x"C3",x"D1",x"C2",x"C3",x"C6",x"00",x"04",x"05",x"06",x"00",x"00",x"C9",x"C2",x"C6",x"C6",x"C6",x"CE",x"BB",x"C2",x"CA",x"C6",x"00",x"05",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"09",x"04",x"0A",x"03",x"00",x"01",x"06",x"00",x"01",x"04",x"00",x"00",x"C6",x"C7",x"C5",x"BF",x"BC",x"CF",x"C1",x"C3",x"CB",x"C2",x"CB",x"C6",x"00",x"08",x"C9",x"C2",x"BB",x"C8",x"C5",x"C8",x"00",x"0B",x"C4",x"BC",x"C4",x"C7",x"CA",x"BF",x"08",x"00",x"00",x"01",x"00",x"06",x"00",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"DC",x"C1",x"03",x"02",x"00",x"02",x"00",x"00",x"05",x"00",x"05",x"0B",x"C3",x"CC",x"DB",x"BC",x"C3",x"C3",x"CA",x"C8",x"BE",x"C8",x"00",x"05",x"02",x"00",x"08",x"05",x"C4",x"BA",x"C8",x"D0",x"AF",x"DF",x"BD",x"C4",x"C4",x"BE",x"10",x"00",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"00",x"00",x"00",x"0C",x"06",x"00",x"03",x"0A",x"0A",x"00",x"00",x"00",x"CD",x"C7",x"CE",x"C5",x"C3",x"CD",x"C2",x"BD",x"C4",x"C4",x"B5",x"C5",x"09",x"0B",x"C4",x"C7",x"C4",x"C9",x"C0",x"C6",x"00",x"00",x"CB",x"BF",x"C6",x"C9",x"C7",x"BB",x"09",x"00",x"00",x"04",x"00",x"09",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"DC",x"C1",x"03",x"02",x"00",x"02",x"00",x"00",x"00",x"00",x"00",x"02",x"04",x"C7",x"BF",x"CF",x"C6",x"C0",x"C9",x"C9",x"CD",x"00",x"00",x"0B",x"00",x"00",x"00",x"02",x"04",x"C7",x"BF",x"CF",x"C6",x"C0",x"C9",x"C9",x"CD",x"00",x"00",x"0B",x"00",x"03",x"C7",x"BF",x"CE",x"C2",x"C3",x"C8",x"09",x"00",x"00",x"04",x"00",x"09",x"00",x"01",x"00",x"00",x"00",x"02",x"04",x"C7",x"BF",x"CF",x"C7",x"C7",x"C7",x"C7",x"C7",x"C7",x"C7",x"C7",x"06",x"0F",x"BC",x"CC",x"C3",x"BC",x"CF",x"C0",x"06",x"0F",x"BC",x"CC",x"C3",x"BC",x"CF",x"C0",x"09",x"00",x"00",x"04",x"00",x"09",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"DC",x"C1",x"03",x"02",x"00",x"02",x"00",x"00",x"00",x"04",x"00",x"00",x"06",x"04",x"16",x"00",x"12",x"00",x"00",x"00",x"07",x"0E",x"00",x"0A",x"00",x"04",x"00",x"00",x"06",x"04",x"16",x"00",x"12",x"00",x"00",x"00",x"07",x"0E",x"00",x"0A",x"00",x"03",x"17",x"00",x"00",x"00",x"02",x"02",x"08",x"00",x"00",x"01",x"00",x"06",x"00",x"04",x"00",x"04",x"00",x"00",x"06",x"04",x"16",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"0A",x"00",x"10",x"03",x"04",x"18",x"00",x"00",x"0A",x"00",x"10",x"03",x"04",x"18",x"08",x"00",x"00",x"01",x"00",x"06",x"00",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"DC",x"C1",x"03",x"02",x"00",x"02",x"00",x"00",x"05",x"0F",x"0D",x"09",x"00",x"00",x"00",x"0E",x"00",x"0D",x"00",x"00",x"00",x"04",x"00",x"00",x"05",x"0F",x"0D",x"09",x"00",x"00",x"00",x"0E",x"00",x"0D",x"00",x"00",x"00",x"04",x"00",x"00",x"00",x"01",x"00",x"0D",x"05",x"00",x"00",x"00",x"00",x"04",x"00",x"02",x"00",x"02",x"00",x"05",x"05",x"0F",x"0D",x"09",x"00",x"00",x"00",x"0E",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"00",x"08",x"00",x"02",x"02",x"00",x"00",x"10",x"00",x"08",x"00",x"02",x"02",x"00",x"00",x"00",x"04",x"00",x"02",x"00",x"02",x"00",x"05",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"DC",x"C1",x"03",x"02",x"00",x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"15",x"05",x"0B",x"00",x"0C",x"00",x"06",x"00",x"0F",x"0D",x"00",x"00",x"00",x"00",x"00",x"00",x"15",x"05",x"0B",x"00",x"0C",x"00",x"06",x"00",x"0F",x"0D",x"00",x"09",x"08",x"00",x"0C",x"05",x"06",x"05",x"00",x"00",x"0C",x"07",x"02",x"00",x"00",x"00",x"06",x"00",x"00",x"00",x"00",x"00",x"15",x"05",x"0B",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"05",x"00",x"00",x"03",x"07",x"02",x"00",x"08",x"05",x"00",x"00",x"03",x"07",x"02",x"00",x"08",x"00",x"0C",x"07",x"02",x"00",x"00",x"00",x"06",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"DC",x"C1",x"03",x"02",x"00",x"02",x"00",x"00",x"00",x"08",x"00",x"00",x"00",x"09",x"04",x"00",x"04",x"0B",x"19",x"00",x"0F",x"00",x"02",x"0A",x"00",x"08",x"00",x"00",x"00",x"09",x"04",x"00",x"04",x"0B",x"19",x"00",x"0F",x"00",x"02",x"0A",x"00",x"08",x"05",x"00",x"00",x"0C",x"13",x"0D",x"00",x"00",x"00",x"03",x"05",x"00",x"00",x"04",x"00",x"08",x"00",x"00",x"00",x"09",x"04",x"00",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"00",x"1D",x"12",x"00",x"00",x"04",x"03",x"0B",x"00",x"1D",x"12",x"00",x"00",x"04",x"03",x"0B",x"00",x"00",x"00",x"03",x"05",x"00",x"00",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"DC",x"C1",x"03",x"02",x"00",x"02",x"00",x"00",x"00",x"00",x"01",x"09",x"0C",x"00",x"16",x"00",x"02",x"04",x"01",x"00",x"00",x"03",x"00",x"16",x"00",x"00",x"01",x"09",x"0C",x"00",x"16",x"00",x"02",x"04",x"01",x"00",x"00",x"03",x"00",x"16",x"00",x"00",x"0C",x"0E",x"00",x"00",x"00",x"00",x"1E",x"14",x"00",x"02",x"02",x"00",x"00",x"0C",x"00",x"00",x"01",x"09",x"0C",x"00",x"16",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"05",x"00",x"00",x"05",x"00",x"03",x"17",x"00",x"05",x"00",x"00",x"05",x"00",x"03",x"17",x"00",x"1E",x"14",x"00",x"02",x"02",x"00",x"00",x"0C",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"DC",x"C1",x"03",x"02",x"00",x"02",x"00",x"00",x"00",x"00",x"0C",x"0C",x"00",x"10",x"00",x"0F",x"00",x"01",x"00",x"01",x"00",x"00",x"20",x"00",x"00",x"00",x"0C",x"0C",x"00",x"10",x"00",x"0F",x"00",x"01",x"00",x"01",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"0B",x"00",x"00",x"0D",x"00",x"02",x"00",x"00",x"07",x"0D",x"00",x"00",x"00",x"00",x"00",x"0C",x"0C",x"00",x"10",x"00",x"0F",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"00",x"00",x"00",x"03",x"06",x"00",x"04",x"00",x"00",x"00",x"00",x"03",x"06",x"00",x"04",x"00",x"02",x"00",x"00",x"07",x"0D",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"DC",x"C1",x"03",x"02",x"00",x"02",x"00",x"00",x"04",x"00",x"03",x"00",x"00",x"00",x"08",x"00",x"00",x"03",x"04",x"08",x"01",x"00",x"00",x"00",x"04",x"00",x"03",x"00",x"00",x"00",x"08",x"00",x"00",x"03",x"04",x"08",x"01",x"00",x"00",x"00",x"04",x"02",x"00",x"04",x"00",x"09",x"0B",x"08",x"00",x"00",x"00",x"01",x"03",x"00",x"00",x"01",x"04",x"00",x"03",x"00",x"00",x"00",x"08",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"06",x"00",x"06",x"00",x"08",x"00",x"11",x"00",x"06",x"00",x"06",x"00",x"08",x"00",x"11",x"00",x"00",x"00",x"00",x"01",x"03",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"DC",x"C1",x"03",x"02",x"00",x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"07",x"05",x"05",x"07",x"00",x"00",x"08",x"09",x"03",x"08",x"00",x"00",x"00",x"17",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"07",x"05",x"00",x"00",x"00",x"17",x"00",x"00",x"00",x"00",x"04",x"00",x"1C",x"09",x"00",x"00",x"03",x"00",x"00",x"00",x"00",x"17",x"00",x"00",x"00",x"00",x"04",x"00",x"1C",x"09",x"00",x"00",x"03",x"00",x"06",x"00",x"0E",x"10",x"00",x"03",x"0C",x"01",x"00",x"00",x"00",x"17",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"00",x"1C",x"09",x"00",x"00",x"03",x"00",x"00",x"00",x"00",x"17",x"00",x"00",x"00",x"00",x"04",x"00",x"1C",x"09",x"00",x"00",x"03",x"00",x"00",x"00",x"00",x"17",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"07",x"05",x"00",x"00",x"00",x"17",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"07",x"05",x"00",x"00",x"00",x"17",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"DC",x"C1",x"03",x"02",x"00",x"02",x"00",x"00",x"00",x"12",x"0D",x"00",x"0D",x"D0",x"C7",x"BA",x"C4",x"BB",x"06",x"03",x"00",x"00",x"01",x"00",x"DE",x"BE",x"BC",x"CD",x"C6",x"00",x"00",x"06",x"00",x"12",x"0D",x"00",x"0D",x"D0",x"C7",x"BA",x"DE",x"BE",x"BC",x"CD",x"C6",x"00",x"00",x"06",x"00",x"08",x"AF",x"B3",x"C3",x"C2",x"CA",x"CC",x"DE",x"BE",x"BC",x"CD",x"C6",x"00",x"00",x"06",x"00",x"08",x"AF",x"B3",x"C3",x"C2",x"CA",x"CC",x"00",x"0C",x"00",x"00",x"00",x"BA",x"BF",x"BE",x"DE",x"BE",x"BC",x"CD",x"C6",x"00",x"00",x"06",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"AF",x"B3",x"C3",x"C2",x"CA",x"CC",x"DE",x"BE",x"BC",x"CD",x"C6",x"00",x"00",x"06",x"00",x"08",x"AF",x"B3",x"C3",x"C2",x"CA",x"CC",x"DE",x"BE",x"BC",x"CD",x"C6",x"00",x"00",x"06",x"00",x"12",x"0D",x"00",x"0D",x"D0",x"C7",x"BA",x"DE",x"BE",x"BC",x"CD",x"C6",x"00",x"00",x"06",x"00",x"12",x"0D",x"00",x"0D",x"D0",x"C7",x"BA",x"DE",x"BE",x"BC",x"CD",x"C6",x"00",x"00",x"06",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"DC",x"C1",x"03",x"02",x"00",x"02",x"00",x"00",x"00",x"00",x"07",x"08",x"C2",x"C8",x"BC",x"CE",x"C7",x"CA",x"C4",x"08",x"00",x"00",x"08",x"CB",x"C4",x"BB",x"C7",x"B1",x"C6",x"CA",x"00",x"05",x"00",x"00",x"07",x"08",x"C2",x"C8",x"BC",x"CE",x"C4",x"BB",x"C7",x"B1",x"C6",x"CA",x"00",x"05",x"00",x"00",x"CB",x"C6",x"CE",x"C5",x"C5",x"BF",x"C4",x"BB",x"C7",x"B1",x"C6",x"CA",x"00",x"05",x"00",x"00",x"CB",x"C6",x"CE",x"C5",x"C5",x"BF",x"02",x"05",x"00",x"01",x"C3",x"D0",x"CD",x"C2",x"C4",x"BB",x"C7",x"B1",x"C6",x"CA",x"00",x"05",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"CB",x"C6",x"CE",x"C5",x"C5",x"BF",x"C4",x"BB",x"C7",x"B1",x"C6",x"CA",x"00",x"05",x"00",x"00",x"CB",x"C6",x"CE",x"C5",x"C5",x"BF",x"C4",x"BB",x"C7",x"B1",x"C6",x"CA",x"00",x"05",x"00",x"00",x"07",x"08",x"C2",x"C8",x"BC",x"CE",x"C4",x"BB",x"C7",x"B1",x"C6",x"CA",x"00",x"05",x"00",x"00",x"07",x"08",x"C2",x"C8",x"BC",x"CE",x"C4",x"BB",x"C7",x"B1",x"C6",x"CA",x"00",x"05",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"DC",x"C1",x"03",x"02",x"00",x"02",x"00",x"00",x"0B",x"06",x"09",x"00",x"BA",x"B0",x"C9",x"B7",x"C7",x"C8",x"C6",x"00",x"00",x"08",x"00",x"D1",x"CF",x"BD",x"C5",x"D2",x"C3",x"CC",x"03",x"07",x"0B",x"06",x"09",x"00",x"BA",x"B0",x"C9",x"B7",x"CF",x"BD",x"C5",x"D2",x"C3",x"CC",x"03",x"07",x"08",x"0A",x"C5",x"CC",x"CD",x"C2",x"C4",x"B5",x"CF",x"BD",x"C5",x"D2",x"C3",x"CC",x"03",x"07",x"08",x"0A",x"C5",x"CC",x"CD",x"C2",x"C4",x"B5",x"00",x"00",x"04",x"00",x"CF",x"C3",x"CF",x"C0",x"CF",x"BD",x"C5",x"D2",x"C3",x"CC",x"03",x"07",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"0A",x"C5",x"CC",x"CD",x"C2",x"C4",x"B5",x"CF",x"BD",x"C5",x"D2",x"C3",x"CC",x"03",x"07",x"08",x"0A",x"C5",x"CC",x"CD",x"C2",x"C4",x"B5",x"CF",x"BD",x"C5",x"D2",x"C3",x"CC",x"03",x"07",x"0B",x"06",x"09",x"00",x"BA",x"B0",x"C9",x"B7",x"CF",x"BD",x"C5",x"D2",x"C3",x"CC",x"03",x"07",x"0B",x"06",x"09",x"00",x"BA",x"B0",x"C9",x"B7",x"CF",x"BD",x"C5",x"D2",x"C3",x"CC",x"03",x"07",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"DC",x"C1",x"03",x"02",x"00",x"02",x"00",x"00",x"00",x"07",x"00",x"C2",x"D1",x"D0",x"BC",x"C7",x"C0",x"D0",x"BF",x"BA",x"0E",x"00",x"CB",x"D0",x"B6",x"D0",x"C3",x"C2",x"D4",x"B8",x"CA",x"05",x"00",x"07",x"00",x"C2",x"D1",x"D0",x"BC",x"C7",x"B6",x"D0",x"C3",x"C2",x"D4",x"B8",x"CA",x"05",x"00",x"0E",x"BC",x"CA",x"CC",x"C4",x"CD",x"C6",x"B6",x"D0",x"C3",x"C2",x"D4",x"B8",x"CA",x"05",x"00",x"0E",x"BC",x"CA",x"CC",x"C4",x"CD",x"C6",x"00",x"00",x"09",x"C8",x"B8",x"D0",x"BA",x"C8",x"B6",x"D0",x"C3",x"C2",x"D4",x"B8",x"CA",x"05",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"0E",x"BC",x"CA",x"CC",x"C4",x"CD",x"C6",x"B6",x"D0",x"C3",x"C2",x"D4",x"B8",x"CA",x"05",x"00",x"0E",x"BC",x"CA",x"CC",x"C4",x"CD",x"C6",x"B6",x"D0",x"C3",x"C2",x"D4",x"B8",x"CA",x"05",x"00",x"07",x"00",x"C2",x"D1",x"D0",x"BC",x"C7",x"B6",x"D0",x"C3",x"C2",x"D4",x"B8",x"CA",x"05",x"00",x"07",x"00",x"C2",x"D1",x"D0",x"BC",x"C7",x"B6",x"D0",x"C3",x"C2",x"D4",x"B8",x"CA",x"05",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"DC",x"C1",x"03",x"02",x"00",x"02",x"00",x"00",x"0C",x"04",x"00",x"D0",x"CF",x"B9",x"C6",x"E1",x"BB",x"C8",x"D1",x"CE",x"0F",x"00",x"B4",x"AF",x"C5",x"D8",x"CC",x"BA",x"B6",x"CE",x"C5",x"00",x"0C",x"04",x"00",x"D0",x"CF",x"B9",x"C6",x"E1",x"C5",x"D8",x"CC",x"BA",x"B6",x"CE",x"C5",x"00",x"00",x"00",x"B4",x"B1",x"C1",x"BE",x"C7",x"CB",x"C5",x"D8",x"CC",x"BA",x"B6",x"CE",x"C5",x"00",x"00",x"00",x"B4",x"B1",x"C1",x"BE",x"C7",x"CB",x"13",x"00",x"00",x"BF",x"C1",x"D9",x"BD",x"C2",x"C5",x"D8",x"CC",x"BA",x"B6",x"CE",x"C5",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"B4",x"B1",x"C1",x"BE",x"C7",x"CB",x"C5",x"D8",x"CC",x"BA",x"B6",x"CE",x"C5",x"00",x"00",x"00",x"B4",x"B1",x"C1",x"BE",x"C7",x"CB",x"C5",x"D8",x"CC",x"BA",x"B6",x"CE",x"C5",x"00",x"0C",x"04",x"00",x"D0",x"CF",x"B9",x"C6",x"E1",x"C5",x"D8",x"CC",x"BA",x"B6",x"CE",x"C5",x"00",x"0C",x"04",x"00",x"D0",x"CF",x"B9",x"C6",x"E1",x"C5",x"D8",x"CC",x"BA",x"B6",x"CE",x"C5",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"DC",x"C1",x"03",x"02",x"00",x"02",x"00",x"00",x"00",x"00",x"B7",x"C2",x"C9",x"BD",x"D1",x"AB",x"C1",x"BC",x"C5",x"C1",x"B5",x"CD",x"C0",x"D3",x"B8",x"BA",x"CA",x"D8",x"BB",x"CA",x"BB",x"D0",x"00",x"00",x"B7",x"C2",x"C9",x"BD",x"D1",x"AB",x"B8",x"BA",x"CA",x"D8",x"BB",x"CA",x"BB",x"D0",x"0A",x"08",x"C2",x"C0",x"CD",x"C4",x"C3",x"BC",x"B8",x"BA",x"CA",x"D8",x"BB",x"CA",x"BB",x"D0",x"0A",x"08",x"C2",x"C0",x"CD",x"C4",x"C3",x"BC",x"0B",x"0C",x"C4",x"CE",x"BD",x"BB",x"CA",x"BD",x"B8",x"BA",x"CA",x"D8",x"BB",x"CA",x"BB",x"D0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"0A",x"08",x"C2",x"C0",x"CD",x"C4",x"C3",x"BC",x"B8",x"BA",x"CA",x"D8",x"BB",x"CA",x"BB",x"D0",x"0A",x"08",x"C2",x"C0",x"CD",x"C4",x"C3",x"BC",x"B8",x"BA",x"CA",x"D8",x"BB",x"CA",x"BB",x"D0",x"00",x"00",x"B7",x"C2",x"C9",x"BD",x"D1",x"AB",x"B8",x"BA",x"CA",x"D8",x"BB",x"CA",x"BB",x"D0",x"00",x"00",x"B7",x"C2",x"C9",x"BD",x"D1",x"AB",x"B8",x"BA",x"CA",x"D8",x"BB",x"CA",x"BB",x"D0",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"DC",x"C1",x"03",x"02",x"00",x"02",x"00",x"00",x"03",x"00",x"D1",x"C7",x"B5",x"D0",x"C3",x"C1",x"D2",x"BD",x"D3",x"C0",x"BD",x"C1",x"C6",x"C7",x"C9",x"CE",x"C5",x"BB",x"D6",x"C6",x"B7",x"CF",x"03",x"00",x"D1",x"C7",x"B5",x"D0",x"C3",x"C1",x"C9",x"CE",x"C5",x"BB",x"D6",x"C6",x"B7",x"CF",x"00",x"05",x"BF",x"CE",x"CC",x"C3",x"CA",x"BC",x"C9",x"CE",x"C5",x"BB",x"D6",x"C6",x"B7",x"CF",x"00",x"05",x"BF",x"CE",x"CC",x"C3",x"CA",x"BC",x"00",x"03",x"BC",x"CA",x"C5",x"D6",x"B5",x"CE",x"C9",x"CE",x"C5",x"BB",x"D6",x"C6",x"B7",x"CF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"05",x"BF",x"CE",x"CC",x"C3",x"CA",x"BC",x"C9",x"CE",x"C5",x"BB",x"D6",x"C6",x"B7",x"CF",x"00",x"05",x"BF",x"CE",x"CC",x"C3",x"CA",x"BC",x"C9",x"CE",x"C5",x"BB",x"D6",x"C6",x"B7",x"CF",x"03",x"00",x"D1",x"C7",x"B5",x"D0",x"C3",x"C1",x"C9",x"CE",x"C5",x"BB",x"D6",x"C6",x"B7",x"CF",x"03",x"00",x"D1",x"C7",x"B5",x"D0",x"C3",x"C1",x"C9",x"CE",x"C5",x"BB",x"D6",x"C6",x"B7",x"CF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"DC",x"C1",x"03",x"02",x"00",x"02",x"00",x"00",x"00",x"00",x"C7",x"C3",x"C4",x"C9",x"BF",x"C8",x"C9",x"C3",x"C3",x"CA",x"B2",x"D6",x"C2",x"CB",x"C9",x"C3",x"C3",x"CA",x"B2",x"D6",x"C2",x"CB",x"2D",x"00",x"BF",x"C3",x"C7",x"C6",x"C6",x"C8",x"C9",x"C3",x"C3",x"CA",x"B2",x"D6",x"C2",x"CB",x"2D",x"00",x"BF",x"C3",x"C7",x"C6",x"C6",x"C8",x"C9",x"C3",x"C3",x"CA",x"B2",x"D6",x"C2",x"CB",x"2D",x"00",x"BF",x"C3",x"C7",x"C6",x"C6",x"C8",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"C9",x"C3",x"C3",x"CA",x"B2",x"D6",x"C2",x"CB",x"2C",x"00",x"00",x"03",x"00",x"00",x"02",x"02",x"00",x"00",x"C7",x"C3",x"C4",x"C9",x"BF",x"C8",x"C9",x"C3",x"C3",x"CA",x"B2",x"D6",x"C2",x"CB",x"2D",x"00",x"BF",x"C3",x"C7",x"C6",x"C6",x"C8",x"C9",x"C3",x"C3",x"CA",x"B2",x"D6",x"C2",x"CB",x"2D",x"00",x"BF",x"C3",x"C7",x"C6",x"C6",x"C8",x"C9",x"C3",x"C3",x"CA",x"B2",x"D6",x"C2",x"CB",x"2D",x"00",x"BF",x"C3",x"C7",x"C6",x"C6",x"C8",x"C9",x"C3",x"C3",x"CA",x"B2",x"D6",x"C2",x"CB",x"2C",x"00",x"00",x"03",x"00",x"00",x"02",x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"DC",x"C1",x"03",x"02",x"00",x"02",x"00",x"00",x"00",x"00",x"C7",x"C3",x"C4",x"C9",x"BF",x"C8",x"00",x"00",x"CD",x"CE",x"B6",x"CB",x"C2",x"C0",x"00",x"00",x"CD",x"CE",x"B6",x"CB",x"C2",x"C0",x"00",x"00",x"CD",x"C4",x"C4",x"C7",x"C7",x"C1",x"00",x"00",x"CD",x"CE",x"B6",x"CB",x"C2",x"C0",x"00",x"00",x"CD",x"C4",x"C4",x"C7",x"C7",x"C1",x"00",x"00",x"CD",x"CE",x"B6",x"CB",x"C2",x"C0",x"00",x"00",x"CD",x"C4",x"C4",x"C7",x"C7",x"C1",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"00",x"00",x"CD",x"CE",x"B6",x"CB",x"C2",x"C0",x"00",x"00",x"06",x"02",x"00",x"01",x"02",x"00",x"00",x"00",x"C7",x"C3",x"C4",x"C9",x"BF",x"C8",x"00",x"00",x"CD",x"CE",x"B6",x"CB",x"C2",x"C0",x"00",x"00",x"CD",x"C4",x"C4",x"C7",x"C7",x"C1",x"00",x"00",x"CD",x"CE",x"B6",x"CB",x"C2",x"C0",x"00",x"00",x"CD",x"C4",x"C4",x"C7",x"C7",x"C1",x"00",x"00",x"CD",x"CE",x"B6",x"CB",x"C2",x"C0",x"00",x"00",x"CD",x"C4",x"C4",x"C7",x"C7",x"C1",x"00",x"00",x"CD",x"CE",x"B6",x"CB",x"C2",x"C0",x"00",x"00",x"06",x"02",x"00",x"01",x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"DC",x"C1",x"03",x"02",x"00",x"02",x"00",x"00",x"00",x"00",x"C7",x"C3",x"C4",x"C9",x"BF",x"C8",x"07",x"0C",x"C6",x"D0",x"C2",x"C1",x"C1",x"CB",x"07",x"0C",x"C6",x"D0",x"C2",x"C1",x"C1",x"CB",x"00",x"07",x"D6",x"C3",x"C5",x"C1",x"C4",x"C7",x"07",x"0C",x"C6",x"D0",x"C2",x"C1",x"C1",x"CB",x"00",x"07",x"D6",x"C3",x"C5",x"C1",x"C4",x"C7",x"07",x"0C",x"C6",x"D0",x"C2",x"C1",x"C1",x"CB",x"00",x"07",x"D6",x"C3",x"C5",x"C1",x"C4",x"C7",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"07",x"0C",x"C6",x"D0",x"C2",x"C1",x"C1",x"CB",x"00",x"09",x"0F",x"00",x"00",x"00",x"00",x"02",x"00",x"00",x"C7",x"C3",x"C4",x"C9",x"BF",x"C8",x"07",x"0C",x"C6",x"D0",x"C2",x"C1",x"C1",x"CB",x"00",x"07",x"D6",x"C3",x"C5",x"C1",x"C4",x"C7",x"07",x"0C",x"C6",x"D0",x"C2",x"C1",x"C1",x"CB",x"00",x"07",x"D6",x"C3",x"C5",x"C1",x"C4",x"C7",x"07",x"0C",x"C6",x"D0",x"C2",x"C1",x"C1",x"CB",x"00",x"07",x"D6",x"C3",x"C5",x"C1",x"C4",x"C7",x"07",x"0C",x"C6",x"D0",x"C2",x"C1",x"C1",x"CB",x"00",x"09",x"0F",x"00",x"00",x"00",x"00",x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"DC",x"C1",x"03",x"02",x"00",x"02",x"00",x"00",x"00",x"00",x"C7",x"C3",x"C4",x"C9",x"BF",x"C8",x"07",x"02",x"C0",x"C9",x"CC",x"BE",x"C1",x"C5",x"07",x"02",x"C0",x"C9",x"CC",x"BE",x"C1",x"C5",x"05",x"0B",x"CD",x"C3",x"CD",x"C0",x"C5",x"C8",x"07",x"02",x"C0",x"C9",x"CC",x"BE",x"C1",x"C5",x"05",x"0B",x"CD",x"C3",x"CD",x"C0",x"C5",x"C8",x"07",x"02",x"C0",x"C9",x"CC",x"BE",x"C1",x"C5",x"05",x"0B",x"CD",x"C3",x"CD",x"C0",x"C5",x"C8",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"07",x"02",x"C0",x"C9",x"CC",x"BE",x"C1",x"C5",x"04",x"0C",x"06",x"01",x"06",x"00",x"00",x"02",x"00",x"00",x"C7",x"C3",x"C4",x"C9",x"BF",x"C8",x"07",x"02",x"C0",x"C9",x"CC",x"BE",x"C1",x"C5",x"05",x"0B",x"CD",x"C3",x"CD",x"C0",x"C5",x"C8",x"07",x"02",x"C0",x"C9",x"CC",x"BE",x"C1",x"C5",x"05",x"0B",x"CD",x"C3",x"CD",x"C0",x"C5",x"C8",x"07",x"02",x"C0",x"C9",x"CC",x"BE",x"C1",x"C5",x"05",x"0B",x"CD",x"C3",x"CD",x"C0",x"C5",x"C8",x"07",x"02",x"C0",x"C9",x"CC",x"BE",x"C1",x"C5",x"04",x"0C",x"06",x"01",x"06",x"00",x"00",x"02",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"DC",x"C1",x"03",x"02",x"00",x"02",x"00",x"00",x"00",x"00",x"C7",x"C3",x"C4",x"C9",x"BF",x"C8",x"02",x"00",x"C0",x"BA",x"CA",x"BF",x"C4",x"C7",x"02",x"00",x"C0",x"BA",x"CA",x"BF",x"C4",x"C7",x"00",x"02",x"C8",x"BF",x"C4",x"C4",x"CE",x"C4",x"02",x"00",x"C0",x"BA",x"CA",x"BF",x"C4",x"C7",x"00",x"02",x"C8",x"BF",x"C4",x"C4",x"CE",x"C4",x"02",x"00",x"C0",x"BA",x"CA",x"BF",x"C4",x"C7",x"00",x"02",x"C8",x"BF",x"C4",x"C4",x"CE",x"C4",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C0",x"BA",x"CA",x"BF",x"C4",x"C7",x"00",x"04",x"02",x"00",x"00",x"00",x"0B",x"00",x"00",x"00",x"C7",x"C3",x"C4",x"C9",x"BF",x"C8",x"02",x"00",x"C0",x"BA",x"CA",x"BF",x"C4",x"C7",x"00",x"02",x"C8",x"BF",x"C4",x"C4",x"CE",x"C4",x"02",x"00",x"C0",x"BA",x"CA",x"BF",x"C4",x"C7",x"00",x"02",x"C8",x"BF",x"C4",x"C4",x"CE",x"C4",x"02",x"00",x"C0",x"BA",x"CA",x"BF",x"C4",x"C7",x"00",x"02",x"C8",x"BF",x"C4",x"C4",x"CE",x"C4",x"02",x"00",x"C0",x"BA",x"CA",x"BF",x"C4",x"C7",x"00",x"04",x"02",x"00",x"00",x"00",x"0B",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"DC",x"C1",x"03",x"02",x"00",x"02",x"00",x"00",x"00",x"00",x"C7",x"C3",x"C4",x"C9",x"BF",x"C8",x"00",x"25",x"AE",x"BE",x"CC",x"CB",x"C4",x"C8",x"00",x"25",x"AE",x"BE",x"CC",x"CB",x"C4",x"C8",x"00",x"01",x"C6",x"BC",x"BF",x"C4",x"D3",x"C4",x"00",x"25",x"AE",x"BE",x"CC",x"CB",x"C4",x"C8",x"00",x"01",x"C6",x"BC",x"BF",x"C4",x"D3",x"C4",x"00",x"25",x"AE",x"BE",x"CC",x"CB",x"C4",x"C8",x"00",x"01",x"C6",x"BC",x"BF",x"C4",x"D3",x"C4",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"00",x"25",x"AE",x"BE",x"CC",x"CB",x"C4",x"C8",x"00",x"03",x"00",x"00",x"00",x"00",x"0F",x"00",x"00",x"00",x"C7",x"C3",x"C4",x"C9",x"BF",x"C8",x"00",x"25",x"AE",x"BE",x"CC",x"CB",x"C4",x"C8",x"00",x"01",x"C6",x"BC",x"BF",x"C4",x"D3",x"C4",x"00",x"25",x"AE",x"BE",x"CC",x"CB",x"C4",x"C8",x"00",x"01",x"C6",x"BC",x"BF",x"C4",x"D3",x"C4",x"00",x"25",x"AE",x"BE",x"CC",x"CB",x"C4",x"C8",x"00",x"01",x"C6",x"BC",x"BF",x"C4",x"D3",x"C4",x"00",x"25",x"AE",x"BE",x"CC",x"CB",x"C4",x"C8",x"00",x"03",x"00",x"00",x"00",x"00",x"0F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"DC",x"C1",x"03",x"02",x"00",x"02",x"00",x"00",x"00",x"00",x"C7",x"C3",x"C4",x"C9",x"BF",x"C8",x"00",x"11",x"C2",x"C2",x"C1",x"C7",x"C4",x"C5",x"00",x"11",x"C2",x"C2",x"C1",x"C7",x"C4",x"C5",x"00",x"00",x"C1",x"BF",x"CC",x"C9",x"C8",x"BD",x"00",x"11",x"C2",x"C2",x"C1",x"C7",x"C4",x"C5",x"00",x"00",x"C1",x"BF",x"CC",x"C9",x"C8",x"BD",x"00",x"11",x"C2",x"C2",x"C1",x"C7",x"C4",x"C5",x"00",x"00",x"C1",x"BF",x"CC",x"C9",x"C8",x"BD",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"00",x"11",x"C2",x"C2",x"C1",x"C7",x"C4",x"C5",x"00",x"00",x"00",x"00",x"06",x"03",x"03",x"00",x"00",x"00",x"C7",x"C3",x"C4",x"C9",x"BF",x"C8",x"00",x"11",x"C2",x"C2",x"C1",x"C7",x"C4",x"C5",x"00",x"00",x"C1",x"BF",x"CC",x"C9",x"C8",x"BD",x"00",x"11",x"C2",x"C2",x"C1",x"C7",x"C4",x"C5",x"00",x"00",x"C1",x"BF",x"CC",x"C9",x"C8",x"BD",x"00",x"11",x"C2",x"C2",x"C1",x"C7",x"C4",x"C5",x"00",x"00",x"C1",x"BF",x"CC",x"C9",x"C8",x"BD",x"00",x"11",x"C2",x"C2",x"C1",x"C7",x"C4",x"C5",x"00",x"00",x"00",x"00",x"06",x"03",x"03",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"DC",x"C1",x"03",x"02",x"00",x"02",x"00",x"00",x"00",x"00",x"C7",x"C3",x"C4",x"C9",x"BF",x"C8",x"06",x"00",x"C7",x"C8",x"CA",x"D5",x"C2",x"BF",x"06",x"00",x"C7",x"C8",x"CA",x"D5",x"C2",x"BF",x"01",x"04",x"CB",x"BD",x"CB",x"C7",x"C3",x"BF",x"06",x"00",x"C7",x"C8",x"CA",x"D5",x"C2",x"BF",x"01",x"04",x"CB",x"BD",x"CB",x"C7",x"C3",x"BF",x"06",x"00",x"C7",x"C8",x"CA",x"D5",x"C2",x"BF",x"01",x"04",x"CB",x"BD",x"CB",x"C7",x"C3",x"BF",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"06",x"00",x"C7",x"C8",x"CA",x"D5",x"C2",x"BF",x"02",x"07",x"05",x"00",x"04",x"01",x"00",x"00",x"00",x"00",x"C7",x"C3",x"C4",x"C9",x"BF",x"C8",x"06",x"00",x"C7",x"C8",x"CA",x"D5",x"C2",x"BF",x"01",x"04",x"CB",x"BD",x"CB",x"C7",x"C3",x"BF",x"06",x"00",x"C7",x"C8",x"CA",x"D5",x"C2",x"BF",x"01",x"04",x"CB",x"BD",x"CB",x"C7",x"C3",x"BF",x"06",x"00",x"C7",x"C8",x"CA",x"D5",x"C2",x"BF",x"01",x"04",x"CB",x"BD",x"CB",x"C7",x"C3",x"BF",x"06",x"00",x"C7",x"C8",x"CA",x"D5",x"C2",x"BF",x"02",x"07",x"05",x"00",x"04",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"DC",x"C1",x"03",x"02",x"00",x"02",x"00",x"00",x"00",x"00",x"C7",x"C3",x"C4",x"C9",x"BF",x"C8",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"00",x"1E",x"C1",x"CE",x"BC",x"C4",x"D0",x"BE",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"00",x"00",x"05",x"00",x"02",x"02",x"00",x"00",x"C7",x"C3",x"C4",x"C9",x"BF",x"C8",x"00",x"1E",x"C1",x"CE",x"BC",x"C4",x"D0",x"BE",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"00",x"1E",x"C1",x"CE",x"BC",x"C4",x"D0",x"BE",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"05",x"00",x"CA",x"DE",x"B5",x"D0",x"C8",x"BA",x"09",x"00",x"CA",x"C6",x"CD",x"CC",x"B7",x"C8",x"09",x"00",x"00",x"04",x"00",x"09",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"DC",x"C1",x"03",x"02",x"00",x"02",x"00",x"00",x"00",x"00",x"C7",x"C3",x"C4",x"C9",x"BF",x"C8",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"00",x"AE",x"C4",x"D1",x"BB",x"C8",x"C7",x"C0",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"00",x"00",x"05",x"00",x"02",x"02",x"00",x"00",x"C7",x"C3",x"C4",x"C9",x"BF",x"C8",x"00",x"AE",x"C4",x"D1",x"BB",x"C8",x"C7",x"C0",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"00",x"AE",x"C4",x"D1",x"BB",x"C8",x"C7",x"C0",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"00",x"00",x"D3",x"BC",x"C8",x"B1",x"D2",x"C7",x"BE",x"07",x"00",x"00",x"0D",x"00",x"00",x"0B",x"08",x"00",x"00",x"01",x"00",x"06",x"00",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"DC",x"C1",x"03",x"02",x"00",x"02",x"00",x"00",x"00",x"00",x"C7",x"C3",x"C4",x"C9",x"BF",x"C8",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"0E",x"B2",x"C9",x"C8",x"BD",x"C3",x"BF",x"C5",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"00",x"00",x"05",x"00",x"02",x"02",x"00",x"00",x"C7",x"C3",x"C4",x"C9",x"BF",x"C8",x"0E",x"B2",x"C9",x"C8",x"BD",x"C3",x"BF",x"C5",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"0E",x"B2",x"C9",x"C8",x"BD",x"C3",x"BF",x"C5",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"00",x"10",x"B9",x"BD",x"C7",x"B6",x"CC",x"C1",x"CB",x"C0",x"03",x"02",x"05",x"00",x"00",x"02",x"00",x"04",x"00",x"02",x"00",x"02",x"00",x"05",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"DC",x"C1",x"03",x"02",x"00",x"02",x"00",x"00",x"00",x"00",x"C7",x"C3",x"C4",x"C9",x"BF",x"C8",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"0C",x"C8",x"C8",x"C6",x"BD",x"C5",x"CC",x"CC",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"00",x"00",x"05",x"00",x"02",x"02",x"00",x"00",x"C7",x"C3",x"C4",x"C9",x"BF",x"C8",x"0C",x"C8",x"C8",x"C6",x"BD",x"C5",x"CC",x"CC",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"0C",x"C8",x"C8",x"C6",x"BD",x"C5",x"CC",x"CC",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"03",x"0E",x"04",x"D3",x"BA",x"C7",x"BE",x"C5",x"D0",x"D4",x"B5",x"B5",x"00",x"00",x"0C",x"11",x"00",x"0C",x"07",x"02",x"00",x"00",x"00",x"06",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"DC",x"C1",x"03",x"02",x"00",x"02",x"00",x"00",x"00",x"00",x"C7",x"C3",x"C4",x"C9",x"BF",x"C8",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"10",x"BA",x"C7",x"CE",x"BA",x"C7",x"CA",x"00",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"00",x"00",x"05",x"00",x"02",x"02",x"00",x"00",x"C7",x"C3",x"C4",x"C9",x"BF",x"C8",x"10",x"BA",x"C7",x"CE",x"BA",x"C7",x"CA",x"00",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"10",x"BA",x"C7",x"CE",x"BA",x"C7",x"CA",x"00",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"15",x"04",x"00",x"C9",x"CD",x"B9",x"CE",x"CC",x"C5",x"B8",x"D6",x"B7",x"D5",x"D1",x"04",x"00",x"00",x"00",x"00",x"03",x"05",x"00",x"00",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"DC",x"C1",x"03",x"02",x"00",x"02",x"00",x"00",x"00",x"00",x"C7",x"C3",x"C4",x"C9",x"BF",x"C8",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"03",x"C4",x"BD",x"C2",x"C4",x"CE",x"00",x"00",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"00",x"00",x"05",x"00",x"02",x"02",x"00",x"00",x"C7",x"C3",x"C4",x"C9",x"BF",x"C8",x"03",x"C4",x"BD",x"C2",x"C4",x"CE",x"00",x"00",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"03",x"C4",x"BD",x"C2",x"C4",x"CE",x"00",x"00",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"00",x"00",x"00",x"15",x"CE",x"CA",x"B8",x"C2",x"CC",x"BD",x"C6",x"CB",x"BF",x"CC",x"BC",x"01",x"1E",x"14",x"00",x"02",x"02",x"00",x"00",x"0C",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"DC",x"C1",x"03",x"02",x"00",x"02",x"00",x"00",x"00",x"00",x"C7",x"C3",x"C4",x"C9",x"BF",x"C8",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"00",x"C8",x"C2",x"C5",x"C6",x"C6",x"C2",x"00",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"00",x"00",x"05",x"00",x"02",x"02",x"00",x"00",x"C7",x"C3",x"C4",x"C9",x"BF",x"C8",x"00",x"C8",x"C2",x"C5",x"C6",x"C6",x"C2",x"00",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"00",x"C8",x"C2",x"C5",x"C6",x"C6",x"C2",x"00",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"00",x"00",x"00",x"04",x"00",x"05",x"C6",x"C7",x"B8",x"C7",x"C4",x"CB",x"B7",x"D1",x"C0",x"05",x"02",x"00",x"00",x"07",x"0D",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"DC",x"C1",x"03",x"02",x"00",x"02",x"00",x"00",x"00",x"00",x"C7",x"C3",x"C4",x"C9",x"BF",x"C8",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"07",x"C5",x"C7",x"C2",x"C9",x"C9",x"BA",x"CD",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"00",x"00",x"05",x"00",x"02",x"02",x"00",x"00",x"C7",x"C3",x"C4",x"C9",x"BF",x"C8",x"07",x"C5",x"C7",x"C2",x"C9",x"C9",x"BA",x"CD",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"07",x"C5",x"C7",x"C2",x"C9",x"C9",x"BA",x"CD",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"13",x"0A",x"00",x"08",x"00",x"00",x"04",x"00",x"D5",x"B8",x"C7",x"D1",x"C2",x"C3",x"BF",x"CC",x"00",x"00",x"00",x"01",x"03",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"DC",x"C1",x"03",x"02",x"00",x"02",x"00",x"00",x"00",x"00",x"C7",x"C3",x"C4",x"C9",x"BF",x"C8",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"00",x"29",x"C8",x"CC",x"AE",x"C7",x"CC",x"C1",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"15",x"98",x"D4",x"C4",x"C9",x"C7",x"C0",x"BF",x"00",x"00",x"BE",x"C7",x"C8",x"C2",x"C4",x"C6",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"00",x"00",x"05",x"00",x"02",x"02",x"00",x"00",x"C7",x"C3",x"C4",x"C9",x"BF",x"C8",x"06",x"BE",x"C7",x"CE",x"BD",x"CA",x"BB",x"BE",x"00",x"00",x"BE",x"C7",x"C8",x"C2",x"C4",x"C6",x"15",x"98",x"D4",x"C4",x"C9",x"C7",x"C0",x"BF",x"00",x"00",x"BE",x"C7",x"C8",x"C2",x"C4",x"C6",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"05",x"00",x"02",x"00",x"04",x"12",x"00",x"06",x"00",x"0E",x"C6",x"BD",x"D2",x"C4",x"CE",x"C4",x"00",x"00",x"00",x"01",x"03",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"DC",x"C1",x"03",x"02",x"00",x"02",x"00",x"00",x"00",x"00",x"C7",x"C3",x"C4",x"C9",x"BF",x"C8",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"CA",x"A5",x"D0",x"C3",x"BB",x"CC",x"C5",x"C4",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"07",x"10",x"D2",x"BF",x"C4",x"C8",x"C5",x"C5",x"03",x"00",x"B9",x"CC",x"D0",x"C1",x"BF",x"C5",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"00",x"00",x"05",x"00",x"02",x"02",x"00",x"00",x"C7",x"C3",x"C4",x"C9",x"BF",x"C8",x"05",x"00",x"C5",x"CD",x"C6",x"C5",x"C5",x"C1",x"03",x"00",x"B9",x"CC",x"D0",x"C1",x"BF",x"C5",x"07",x"10",x"D2",x"BF",x"C4",x"C8",x"C5",x"C5",x"03",x"00",x"B9",x"CC",x"D0",x"C1",x"BF",x"C5",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"00",x"0D",x"BE",x"B5",x"C5",x"BA",x"BF",x"DA",x"08",x"12",x"C3",x"AE",x"C7",x"D4",x"B1",x"C9",x"02",x"00",x"00",x"07",x"0D",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"DC",x"C1",x"03",x"02",x"00",x"02",x"00",x"00",x"00",x"00",x"C7",x"C3",x"C4",x"C9",x"BF",x"C8",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"C9",x"BA",x"C9",x"C3",x"C3",x"C9",x"C0",x"C8",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"01",x"00",x"CA",x"C1",x"BF",x"CC",x"C5",x"C7",x"1F",x"18",x"C1",x"C7",x"C6",x"B9",x"C1",x"D1",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"00",x"00",x"05",x"00",x"02",x"02",x"00",x"00",x"C7",x"C3",x"C4",x"C9",x"BF",x"C8",x"07",x"02",x"C9",x"C0",x"C6",x"CB",x"C8",x"C4",x"1F",x"18",x"C1",x"C7",x"C6",x"B9",x"C1",x"D1",x"01",x"00",x"CA",x"C1",x"BF",x"CC",x"C5",x"C7",x"1F",x"18",x"C1",x"C7",x"C6",x"B9",x"C1",x"D1",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"04",x"00",x"DC",x"D0",x"C6",x"B9",x"BF",x"C4",x"00",x"00",x"B0",x"CC",x"C3",x"BC",x"BE",x"C8",x"1E",x"14",x"00",x"02",x"02",x"00",x"00",x"0C",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"DC",x"C1",x"03",x"02",x"00",x"02",x"00",x"00",x"00",x"00",x"C7",x"C3",x"C4",x"C9",x"BF",x"C8",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"BF",x"D1",x"CB",x"C0",x"C2",x"C6",x"BF",x"CA",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"00",x"07",x"BD",x"BF",x"BD",x"CD",x"C6",x"C7",x"00",x"00",x"BD",x"C8",x"C8",x"C2",x"C4",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"00",x"00",x"05",x"00",x"02",x"02",x"00",x"00",x"C7",x"C3",x"C4",x"C9",x"BF",x"C8",x"02",x"02",x"CE",x"B5",x"CD",x"C9",x"C9",x"C4",x"00",x"00",x"BD",x"C8",x"C8",x"C2",x"C4",x"C9",x"00",x"07",x"BD",x"BF",x"BD",x"CD",x"C6",x"C7",x"00",x"00",x"BD",x"C8",x"C8",x"C2",x"C4",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"09",x"00",x"C3",x"D2",x"C8",x"C7",x"CF",x"BD",x"01",x"10",x"C4",x"C8",x"D1",x"CC",x"C2",x"C5",x"00",x"00",x"00",x"03",x"05",x"00",x"00",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"DC",x"C1",x"03",x"02",x"00",x"02",x"00",x"00",x"00",x"00",x"C7",x"C3",x"C4",x"C9",x"BF",x"C8",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"BF",x"D2",x"BB",x"C4",x"D2",x"C8",x"BB",x"C8",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"00",x"00",x"C8",x"C1",x"C7",x"C8",x"C7",x"C3",x"00",x"12",x"C8",x"C7",x"C1",x"C2",x"C4",x"CB",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"00",x"00",x"05",x"00",x"02",x"02",x"00",x"00",x"C7",x"C3",x"C4",x"C9",x"BF",x"C8",x"00",x"00",x"C5",x"B5",x"CC",x"BE",x"CB",x"BF",x"00",x"12",x"C8",x"C7",x"C1",x"C2",x"C4",x"CB",x"00",x"00",x"C8",x"C1",x"C7",x"C8",x"C7",x"C3",x"00",x"12",x"C8",x"C7",x"C1",x"C2",x"C4",x"CB",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"00",x"00",x"C0",x"C7",x"C6",x"BA",x"CE",x"C9",x"00",x"00",x"BF",x"C8",x"C1",x"CA",x"D4",x"C2",x"00",x"0C",x"07",x"02",x"00",x"00",x"00",x"06",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"DC",x"C1",x"03",x"02",x"00",x"02",x"00",x"00",x"00",x"00",x"C7",x"C3",x"C4",x"C9",x"BF",x"C8",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"C5",x"D7",x"BB",x"C5",x"CC",x"C1",x"C0",x"CC",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"05",x"06",x"D0",x"C2",x"C9",x"C5",x"C7",x"BE",x"00",x"08",x"C1",x"C8",x"C2",x"C5",x"BF",x"CA",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"00",x"00",x"05",x"00",x"02",x"02",x"00",x"00",x"C7",x"C3",x"C4",x"C9",x"BF",x"C8",x"00",x"23",x"C7",x"B6",x"C5",x"BD",x"C6",x"C0",x"00",x"08",x"C1",x"C8",x"C2",x"C5",x"BF",x"CA",x"05",x"06",x"D0",x"C2",x"C9",x"C5",x"C7",x"BE",x"00",x"08",x"C1",x"C8",x"C2",x"C5",x"BF",x"CA",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"08",x"04",x"C3",x"B9",x"BE",x"B7",x"BF",x"CB",x"00",x"0E",x"C1",x"CF",x"C1",x"BA",x"C3",x"C4",x"00",x"04",x"00",x"02",x"00",x"02",x"00",x"05",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"DC",x"C1",x"03",x"02",x"00",x"02",x"00",x"00",x"00",x"00",x"C7",x"C3",x"C4",x"C9",x"BF",x"C8",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"BB",x"CE",x"BB",x"C5",x"CA",x"C5",x"C8",x"C0",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"00",x"0B",x"C4",x"BC",x"C4",x"C7",x"CA",x"BF",x"09",x"00",x"BA",x"C7",x"C3",x"C9",x"B9",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"00",x"00",x"05",x"00",x"02",x"02",x"00",x"00",x"C7",x"C3",x"C4",x"C9",x"BF",x"C8",x"00",x"02",x"CF",x"C2",x"CB",x"BE",x"BE",x"CA",x"09",x"00",x"BA",x"C7",x"C3",x"C9",x"B9",x"C9",x"00",x"0B",x"C4",x"BC",x"C4",x"C7",x"CA",x"BF",x"09",x"00",x"BA",x"C7",x"C3",x"C9",x"B9",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"0C",x"00",x"BE",x"C4",x"C5",x"C7",x"BC",x"BD",x"09",x"0D",x"C9",x"BB",x"B7",x"C8",x"C6",x"C3",x"08",x"00",x"00",x"01",x"00",x"06",x"00",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"DC",x"C1",x"03",x"02",x"00",x"02",x"00",x"00",x"00",x"00",x"C7",x"C3",x"C4",x"C9",x"BF",x"C8",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"C1",x"CB",x"BC",x"C6",x"C6",x"BF",x"CD",x"C6",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"00",x"00",x"CB",x"BF",x"C6",x"C9",x"C7",x"BB",x"0A",x"00",x"BC",x"C8",x"C1",x"CB",x"B9",x"C6",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"00",x"00",x"05",x"00",x"02",x"02",x"00",x"00",x"C7",x"C3",x"C4",x"C9",x"BF",x"C8",x"07",x"00",x"C2",x"D0",x"C9",x"C2",x"C1",x"C8",x"0A",x"00",x"BC",x"C8",x"C1",x"CB",x"B9",x"C6",x"00",x"00",x"CB",x"BF",x"C6",x"C9",x"C7",x"BB",x"0A",x"00",x"BC",x"C8",x"C1",x"CB",x"B9",x"C6",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"00",x"00",x"C6",x"CD",x"CE",x"C1",x"D0",x"C0",x"00",x"06",x"C5",x"CA",x"CA",x"B4",x"DB",x"C3",x"09",x"00",x"00",x"04",x"00",x"09",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
		(x"DC",x"C1",x"03",x"02",x"00",x"02",x"00",x"00",x"00",x"00",x"C7",x"C3",x"C4",x"C9",x"BF",x"C8",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"C9",x"C3",x"C3",x"CA",x"B2",x"D6",x"C2",x"CB",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"00",x"02",x"C6",x"C7",x"BF",x"CB",x"B9",x"C9",x"00",x"18",x"C7",x"D1",x"B4",x"CE",x"C3",x"C5",x"02",x"00",x"00",x"00",x"05",x"00",x"02",x"02",x"00",x"00",x"C7",x"C3",x"C4",x"C9",x"BF",x"C8",x"00",x"13",x"C7",x"C2",x"B5",x"D5",x"BE",x"C3",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"00",x"02",x"C6",x"C7",x"BF",x"CB",x"B9",x"C9",x"00",x"18",x"C7",x"D1",x"B4",x"CE",x"C3",x"C5",x"00",x"02",x"C6",x"C7",x"BF",x"CB",x"B9",x"C9",x"00",x"18",x"C7",x"D1",x"B4",x"CE",x"C3",x"C5",x"07",x"00",x"21",x"07",x"00",x"00",x"00",x"07",x"00",x"05",x"02",x"02",x"01",x"00",x"06",x"01"),
		(x"DC",x"C1",x"03",x"02",x"00",x"02",x"00",x"00",x"00",x"00",x"C7",x"C3",x"C4",x"C9",x"BF",x"C8",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"00",x"00",x"CD",x"CE",x"B6",x"CB",x"C2",x"C0",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"05",x"09",x"C0",x"CE",x"C1",x"C6",x"C2",x"CA",x"C4",x"AA",x"C5",x"C3",x"B7",x"D3",x"CE",x"B9",x"02",x"00",x"00",x"00",x"05",x"00",x"02",x"02",x"00",x"00",x"C7",x"C3",x"C4",x"C9",x"BF",x"C8",x"09",x"AB",x"C4",x"C3",x"C3",x"CD",x"BB",x"C4",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"05",x"09",x"C0",x"CE",x"C1",x"C6",x"C2",x"CA",x"C4",x"AA",x"C5",x"C3",x"B7",x"D3",x"CE",x"B9",x"05",x"09",x"C0",x"CE",x"C1",x"C6",x"C2",x"CA",x"C4",x"AA",x"C5",x"C3",x"B7",x"D3",x"CE",x"B9",x"04",x"01",x"B4",x"B2",x"C5",x"C1",x"C5",x"D3",x"00",x"01",x"04",x"03",x"00",x"00",x"04",x"00"),
		(x"DC",x"C1",x"03",x"02",x"00",x"02",x"00",x"00",x"00",x"00",x"C7",x"C3",x"C4",x"C9",x"BF",x"C8",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"07",x"0C",x"C6",x"D0",x"C2",x"C1",x"C1",x"CB",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"04",x"00",x"BA",x"CE",x"C8",x"CB",x"BF",x"CB",x"C6",x"CA",x"C3",x"BE",x"C4",x"CA",x"CA",x"BC",x"02",x"00",x"00",x"00",x"05",x"00",x"02",x"02",x"00",x"00",x"C7",x"C3",x"C4",x"C9",x"BF",x"C8",x"05",x"C6",x"C5",x"CF",x"C4",x"C9",x"C2",x"BF",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"04",x"00",x"BA",x"CE",x"C8",x"CB",x"BF",x"CB",x"C6",x"CA",x"C3",x"BE",x"C4",x"CA",x"CA",x"BC",x"04",x"00",x"BA",x"CE",x"C8",x"CB",x"BF",x"CB",x"C6",x"CA",x"C3",x"BE",x"C4",x"CA",x"CA",x"BC",x"00",x"00",x"CF",x"C4",x"D0",x"C4",x"C1",x"C6",x"06",x"00",x"00",x"04",x"00",x"03",x"00",x"00"),
		(x"DC",x"C1",x"03",x"02",x"00",x"02",x"00",x"00",x"00",x"00",x"C7",x"C3",x"C4",x"C9",x"BF",x"C8",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"07",x"02",x"C0",x"C9",x"CC",x"BE",x"C1",x"C5",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"04",x"09",x"A2",x"C8",x"C9",x"C6",x"C3",x"C1",x"B8",x"D3",x"C6",x"B9",x"C2",x"CF",x"C0",x"C9",x"02",x"00",x"00",x"00",x"05",x"00",x"02",x"02",x"00",x"00",x"C7",x"C3",x"C4",x"C9",x"BF",x"C8",x"06",x"D1",x"C3",x"CC",x"CA",x"C8",x"C4",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"04",x"09",x"A2",x"C8",x"C9",x"C6",x"C3",x"C1",x"B8",x"D3",x"C6",x"B9",x"C2",x"CF",x"C0",x"C9",x"04",x"09",x"A2",x"C8",x"C9",x"C6",x"C3",x"C1",x"B8",x"D3",x"C6",x"B9",x"C2",x"CF",x"C0",x"C9",x"0A",x"04",x"CA",x"CC",x"CD",x"C0",x"C0",x"BA",x"12",x"00",x"00",x"04",x"01",x"07",x"00",x"00"),
		(x"DC",x"C1",x"03",x"02",x"00",x"02",x"00",x"00",x"00",x"00",x"C7",x"C3",x"C4",x"C9",x"BF",x"C8",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C0",x"BA",x"CA",x"BF",x"C4",x"C7",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"00",x"00",x"19",x"C9",x"BE",x"C8",x"B9",x"C7",x"CC",x"CE",x"BD",x"C0",x"CF",x"C1",x"BE",x"00",x"02",x"00",x"00",x"00",x"05",x"00",x"02",x"02",x"00",x"00",x"C7",x"C3",x"C4",x"C9",x"BF",x"C8",x"00",x"BD",x"C9",x"BB",x"C9",x"C9",x"BC",x"00",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"00",x"00",x"19",x"C9",x"BE",x"C8",x"B9",x"C7",x"CC",x"CE",x"BD",x"C0",x"CF",x"C1",x"BE",x"00",x"00",x"00",x"19",x"C9",x"BE",x"C8",x"B9",x"C7",x"CC",x"CE",x"BD",x"C0",x"CF",x"C1",x"BE",x"00",x"07",x"09",x"C2",x"CA",x"CE",x"C3",x"C8",x"CC",x"22",x"01",x"02",x"03",x"00",x"07",x"00",x"00"),
		(x"DC",x"C1",x"03",x"02",x"00",x"02",x"00",x"00",x"00",x"00",x"C7",x"C3",x"C4",x"C9",x"BF",x"C8",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"00",x"25",x"AE",x"BE",x"CC",x"CB",x"C4",x"C8",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"00",x"00",x"0C",x"C2",x"C3",x"CA",x"BC",x"C1",x"C2",x"C5",x"C8",x"C6",x"D2",x"C5",x"BA",x"0D",x"02",x"00",x"00",x"00",x"05",x"00",x"02",x"02",x"00",x"00",x"C7",x"C3",x"C4",x"C9",x"BF",x"C8",x"00",x"BB",x"C5",x"C6",x"BF",x"C8",x"D0",x"04",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"00",x"00",x"0C",x"C2",x"C3",x"CA",x"BC",x"C1",x"C2",x"C5",x"C8",x"C6",x"D2",x"C5",x"BA",x"0D",x"00",x"00",x"0C",x"C2",x"C3",x"CA",x"BC",x"C1",x"C2",x"C5",x"C8",x"C6",x"D2",x"C5",x"BA",x"0D",x"00",x"00",x"B8",x"B1",x"C1",x"BD",x"C3",x"D2",x"00",x"00",x"00",x"04",x"00",x"0F",x"00",x"00"),
		(x"DC",x"C1",x"03",x"02",x"00",x"02",x"00",x"00",x"00",x"00",x"C7",x"C3",x"C4",x"C9",x"BF",x"C8",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"00",x"11",x"C2",x"C2",x"C1",x"C7",x"C4",x"C5",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"05",x"01",x"00",x"00",x"C2",x"CC",x"BD",x"C3",x"C6",x"CE",x"BB",x"C2",x"CA",x"C6",x"00",x"05",x"02",x"00",x"00",x"00",x"05",x"00",x"02",x"02",x"00",x"00",x"C7",x"C3",x"C4",x"C9",x"BF",x"C8",x"05",x"BC",x"C2",x"CC",x"BF",x"C5",x"00",x"02",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"05",x"01",x"00",x"00",x"C2",x"CC",x"BD",x"C3",x"C6",x"CE",x"BB",x"C2",x"CA",x"C6",x"00",x"05",x"05",x"01",x"00",x"00",x"C2",x"CC",x"BD",x"C3",x"C6",x"CE",x"BB",x"C2",x"CA",x"C6",x"00",x"05",x"0C",x"02",x"C8",x"BE",x"CE",x"C2",x"BD",x"C2",x"00",x"05",x"06",x"00",x"00",x"07",x"00",x"03"),
		(x"DC",x"C1",x"03",x"02",x"00",x"02",x"00",x"00",x"00",x"00",x"C7",x"C3",x"C4",x"C9",x"BF",x"C8",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"06",x"00",x"C7",x"C8",x"CA",x"D5",x"C2",x"BF",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"0C",x"00",x"00",x"00",x"CA",x"CD",x"C6",x"C7",x"AF",x"DF",x"BD",x"C4",x"C4",x"BE",x"10",x"00",x"02",x"00",x"00",x"00",x"05",x"00",x"02",x"02",x"00",x"00",x"C7",x"C3",x"C4",x"C9",x"BF",x"C8",x"05",x"C5",x"C6",x"D9",x"BC",x"B6",x"0C",x"00",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"02",x"00",x"C3",x"C3",x"CA",x"C4",x"C1",x"C9",x"0C",x"00",x"00",x"00",x"CA",x"CD",x"C6",x"C7",x"AF",x"DF",x"BD",x"C4",x"C4",x"BE",x"10",x"00",x"0C",x"00",x"00",x"00",x"CA",x"CD",x"C6",x"C7",x"AF",x"DF",x"BD",x"C4",x"C4",x"BE",x"10",x"00",x"00",x"00",x"C5",x"CC",x"CE",x"C0",x"C4",x"C1",x"0C",x"07",x"01",x"05",x"00",x"06",x"00",x"02"),
		(x"D8",x"BD",x"10",x"07",x"00",x"00",x"05",x"01",x"00",x"03",x"C7",x"BF",x"CE",x"C2",x"C3",x"C8",x"06",x"0F",x"BC",x"CC",x"C3",x"BC",x"CF",x"C0",x"06",x"0F",x"BC",x"CC",x"C3",x"BC",x"CF",x"C0",x"06",x"0F",x"BC",x"CC",x"C3",x"BC",x"CF",x"C0",x"06",x"0F",x"BC",x"CC",x"C3",x"BC",x"CF",x"C0",x"06",x"0F",x"BC",x"CC",x"C3",x"BC",x"CF",x"C0",x"06",x"0F",x"BC",x"CC",x"C3",x"BC",x"CF",x"C0",x"06",x"0F",x"BC",x"CC",x"C3",x"BC",x"CF",x"C0",x"07",x"00",x"0C",x"00",x"05",x"C8",x"CC",x"C5",x"C6",x"C0",x"C9",x"C9",x"CD",x"00",x"00",x"0B",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"03",x"C7",x"BF",x"CE",x"C2",x"C3",x"C8",x"00",x"C5",x"D0",x"D2",x"BB",x"02",x"04",x"07",x"00",x"03",x"C7",x"BF",x"CE",x"C2",x"C3",x"C8",x"06",x"0F",x"BC",x"CC",x"C3",x"BC",x"CF",x"C0",x"07",x"00",x"0C",x"00",x"05",x"C8",x"CC",x"C5",x"C6",x"C0",x"C9",x"C9",x"CD",x"00",x"00",x"0B",x"00",x"00",x"00",x"02",x"04",x"C7",x"BF",x"CF",x"C6",x"C0",x"C9",x"C9",x"CD",x"00",x"00",x"0B",x"00",x"03",x"C7",x"BF",x"CE",x"C2",x"C3",x"C8",x"00",x"00",x"01",x"00",x"04",x"10",x"00",x"00"),
		(x"DA",x"BC",x"00",x"16",x"04",x"08",x"00",x"00",x"00",x"03",x"17",x"00",x"00",x"00",x"02",x"02",x"00",x"00",x"0A",x"00",x"10",x"03",x"04",x"18",x"00",x"00",x"0A",x"00",x"10",x"03",x"04",x"18",x"00",x"00",x"0A",x"00",x"10",x"03",x"04",x"18",x"00",x"00",x"0A",x"00",x"10",x"03",x"04",x"18",x"00",x"00",x"0A",x"00",x"10",x"03",x"04",x"18",x"00",x"00",x"0A",x"00",x"10",x"03",x"04",x"18",x"00",x"00",x"0A",x"00",x"10",x"03",x"04",x"18",x"02",x"00",x"0E",x"00",x"0F",x"00",x"00",x"00",x"12",x"00",x"00",x"00",x"07",x"0E",x"00",x"0A",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"03",x"17",x"00",x"00",x"00",x"02",x"02",x"0C",x"00",x"00",x"00",x"05",x"04",x"00",x"04",x"00",x"03",x"17",x"00",x"00",x"00",x"02",x"02",x"00",x"00",x"0A",x"00",x"10",x"03",x"04",x"18",x"02",x"00",x"0E",x"00",x"0F",x"00",x"00",x"00",x"12",x"00",x"00",x"00",x"07",x"0E",x"00",x"0A",x"00",x"04",x"00",x"00",x"06",x"04",x"16",x"00",x"12",x"00",x"00",x"00",x"07",x"0E",x"00",x"0A",x"00",x"03",x"17",x"00",x"00",x"00",x"02",x"02",x"05",x"08",x"0F",x"00",x"04",x"00",x"00",x"06"),
		(x"E9",x"B8",x"08",x"00",x"00",x"05",x"03",x"00",x"00",x"01",x"00",x"0D",x"05",x"00",x"00",x"00",x"10",x"00",x"08",x"00",x"02",x"02",x"00",x"00",x"10",x"00",x"08",x"00",x"02",x"02",x"00",x"00",x"10",x"00",x"08",x"00",x"02",x"02",x"00",x"00",x"10",x"00",x"08",x"00",x"02",x"02",x"00",x"00",x"10",x"00",x"08",x"00",x"02",x"02",x"00",x"00",x"10",x"00",x"08",x"00",x"02",x"02",x"00",x"00",x"10",x"00",x"08",x"00",x"02",x"02",x"00",x"00",x"02",x"01",x"00",x"00",x"01",x"00",x"02",x"09",x"00",x"0D",x"00",x"00",x"00",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"00",x"0D",x"05",x"00",x"00",x"00",x"00",x"00",x"0E",x"00",x"0E",x"0B",x"00",x"01",x"00",x"01",x"00",x"0D",x"05",x"00",x"00",x"00",x"10",x"00",x"08",x"00",x"02",x"02",x"00",x"00",x"02",x"01",x"00",x"00",x"01",x"00",x"02",x"09",x"00",x"0D",x"00",x"00",x"00",x"04",x"00",x"00",x"05",x"0F",x"0D",x"09",x"00",x"00",x"00",x"0E",x"00",x"0D",x"00",x"00",x"00",x"04",x"00",x"00",x"00",x"01",x"00",x"0D",x"05",x"00",x"00",x"00",x"0E",x"07",x"00",x"00",x"06",x"00",x"0A",x"09"),
		(x"DF",x"D6",x"00",x"02",x"02",x"00",x"00",x"06",x"09",x"08",x"00",x"0C",x"05",x"06",x"05",x"00",x"05",x"00",x"00",x"03",x"07",x"02",x"00",x"08",x"05",x"00",x"00",x"03",x"07",x"02",x"00",x"08",x"05",x"00",x"00",x"03",x"07",x"02",x"00",x"08",x"05",x"00",x"00",x"03",x"07",x"02",x"00",x"08",x"05",x"00",x"00",x"03",x"07",x"02",x"00",x"08",x"05",x"00",x"00",x"03",x"07",x"02",x"00",x"08",x"05",x"00",x"00",x"03",x"07",x"02",x"00",x"08",x"00",x"1D",x"08",x"00",x"0A",x"04",x"00",x"0E",x"00",x"0C",x"00",x"06",x"00",x"0F",x"0D",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"09",x"08",x"00",x"0C",x"05",x"06",x"05",x"00",x"04",x"0B",x"04",x"00",x"0B",x"00",x"00",x"0D",x"09",x"08",x"00",x"0C",x"05",x"06",x"05",x"00",x"05",x"00",x"00",x"03",x"07",x"02",x"00",x"08",x"00",x"1D",x"08",x"00",x"0A",x"04",x"00",x"0E",x"00",x"0C",x"00",x"06",x"00",x"0F",x"0D",x"00",x"00",x"00",x"00",x"00",x"00",x"15",x"05",x"0B",x"00",x"0C",x"00",x"06",x"00",x"0F",x"0D",x"00",x"09",x"08",x"00",x"0C",x"05",x"06",x"05",x"00",x"00",x"00",x"00",x"02",x"11",x"08",x"00",x"03"),
		(x"D4",x"CC",x"02",x"04",x"BF",x"BF",x"00",x"09",x"00",x"08",x"05",x"00",x"00",x"0C",x"13",x"0D",x"00",x"1D",x"12",x"00",x"00",x"04",x"03",x"0B",x"00",x"1D",x"12",x"00",x"00",x"04",x"03",x"0B",x"00",x"1D",x"12",x"00",x"00",x"04",x"03",x"0B",x"00",x"1D",x"12",x"00",x"00",x"04",x"03",x"0B",x"00",x"1D",x"12",x"00",x"00",x"04",x"03",x"0B",x"00",x"1D",x"12",x"00",x"00",x"04",x"03",x"0B",x"00",x"1D",x"12",x"00",x"00",x"04",x"03",x"0B",x"0B",x"00",x"00",x"03",x"00",x"0F",x"00",x"00",x"04",x"0B",x"19",x"00",x"0F",x"00",x"02",x"0A",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"08",x"05",x"00",x"00",x"0C",x"13",x"0D",x"04",x"00",x"10",x"00",x"00",x"00",x"00",x"08",x"00",x"08",x"05",x"00",x"00",x"0C",x"13",x"0D",x"00",x"1D",x"12",x"00",x"00",x"04",x"03",x"0B",x"0B",x"00",x"00",x"03",x"00",x"0F",x"00",x"00",x"04",x"0B",x"19",x"00",x"0F",x"00",x"02",x"0A",x"00",x"08",x"00",x"00",x"00",x"09",x"04",x"00",x"04",x"0B",x"19",x"00",x"0F",x"00",x"02",x"0A",x"00",x"08",x"05",x"00",x"00",x"0C",x"13",x"0D",x"01",x"00",x"03",x"00",x"BB",x"BB",x"00",x"0A"),
		(x"D6",x"C4",x"08",x"04",x"BC",x"E4",x"01",x"00",x"00",x"00",x"0C",x"0E",x"00",x"00",x"00",x"00",x"05",x"00",x"00",x"05",x"00",x"03",x"17",x"00",x"05",x"00",x"00",x"05",x"00",x"03",x"17",x"00",x"05",x"00",x"00",x"05",x"00",x"03",x"17",x"00",x"05",x"00",x"00",x"05",x"00",x"03",x"17",x"00",x"05",x"00",x"00",x"05",x"00",x"03",x"17",x"00",x"05",x"00",x"00",x"05",x"00",x"03",x"17",x"00",x"05",x"00",x"00",x"05",x"00",x"03",x"17",x"00",x"03",x"00",x"00",x"02",x"15",x"00",x"0C",x"04",x"02",x"04",x"01",x"00",x"00",x"03",x"00",x"16",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"0C",x"0E",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"07",x"00",x"00",x"0C",x"00",x"00",x"00",x"0C",x"0E",x"00",x"00",x"00",x"00",x"05",x"00",x"00",x"05",x"00",x"03",x"17",x"00",x"03",x"00",x"00",x"02",x"15",x"00",x"0C",x"04",x"02",x"04",x"01",x"00",x"00",x"03",x"00",x"16",x"00",x"00",x"01",x"09",x"0C",x"00",x"16",x"00",x"02",x"04",x"01",x"00",x"00",x"03",x"00",x"16",x"00",x"00",x"0C",x"0E",x"00",x"00",x"00",x"00",x"0E",x"17",x"00",x"15",x"B6",x"B7",x"05",x"01"),
		(x"E5",x"BA",x"0A",x"03",x"00",x"00",x"00",x"02",x"00",x"00",x"00",x"0B",x"00",x"00",x"0D",x"00",x"00",x"00",x"00",x"03",x"06",x"00",x"04",x"00",x"00",x"00",x"00",x"03",x"06",x"00",x"04",x"00",x"00",x"00",x"00",x"03",x"06",x"00",x"04",x"00",x"00",x"00",x"00",x"03",x"06",x"00",x"04",x"00",x"00",x"00",x"00",x"03",x"06",x"00",x"04",x"00",x"00",x"00",x"00",x"03",x"06",x"00",x"04",x"00",x"00",x"00",x"00",x"03",x"06",x"00",x"04",x"00",x"00",x"03",x"0B",x"06",x"00",x"02",x"08",x"00",x"00",x"01",x"00",x"01",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"0B",x"00",x"00",x"0D",x"00",x"05",x"00",x"05",x"10",x"04",x"10",x"00",x"02",x"00",x"00",x"00",x"0B",x"00",x"00",x"0D",x"00",x"00",x"00",x"00",x"03",x"06",x"00",x"04",x"00",x"00",x"03",x"0B",x"06",x"00",x"02",x"08",x"00",x"00",x"01",x"00",x"01",x"00",x"00",x"20",x"00",x"00",x"00",x"0C",x"0C",x"00",x"10",x"00",x"0F",x"00",x"01",x"00",x"01",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"0B",x"00",x"00",x"0D",x"00",x"00",x"00",x"10",x"00",x"0D",x"00",x"01",x"00"),
		(x"DC",x"C3",x"00",x"01",x"0A",x"02",x"00",x"0B",x"04",x"02",x"00",x"04",x"00",x"09",x"0B",x"08",x"06",x"00",x"06",x"00",x"08",x"00",x"11",x"00",x"06",x"00",x"06",x"00",x"08",x"00",x"11",x"00",x"06",x"00",x"06",x"00",x"08",x"00",x"11",x"00",x"06",x"00",x"06",x"00",x"08",x"00",x"11",x"00",x"06",x"00",x"06",x"00",x"08",x"00",x"11",x"00",x"06",x"00",x"06",x"00",x"08",x"00",x"11",x"00",x"06",x"00",x"06",x"00",x"08",x"00",x"11",x"00",x"00",x"05",x"09",x"00",x"00",x"00",x"00",x"07",x"00",x"03",x"04",x"08",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"02",x"00",x"04",x"00",x"09",x"0B",x"08",x"0A",x"06",x"00",x"0B",x"01",x"00",x"03",x"00",x"04",x"02",x"00",x"04",x"00",x"09",x"0B",x"08",x"06",x"00",x"06",x"00",x"08",x"00",x"11",x"00",x"00",x"05",x"09",x"00",x"00",x"00",x"00",x"07",x"00",x"03",x"04",x"08",x"01",x"00",x"00",x"00",x"04",x"00",x"03",x"00",x"00",x"00",x"08",x"00",x"00",x"03",x"04",x"08",x"01",x"00",x"00",x"00",x"04",x"02",x"00",x"04",x"00",x"09",x"0B",x"08",x"03",x"05",x"00",x"00",x"09",x"00",x"00",x"02")
	
	);

begin

	dat_R <= titulo_R( dir_y )( dir_x );
	dat_G <= titulo_G( dir_y )( dir_x );
	dat_B <= titulo_B( dir_y )( dir_x );

end comp;